conectix             1�qemu  Wi2k     `      `     ����u�M���<���                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������                 ���v                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �� |  � �м  h�h 1�1�� ��(  �A��U��r��U�u�� 0�� f1�f1��: �U �$Could not locate active partition
 �� ����t����f`�M r��� �����u�fa�f`&�w&�O&ff�� &��t� r��&�G<t<t<�u��fa� �P� �� r
&�>�U�t�X�� f`1۴���fa�f`�!�%f�>'f�6+��B�fa�                                                                                                                                                                                                             � �?     �  U�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �*� � �м  h�h 1�1�� ��#  �A��U��r��U�u�� � 0�� f1�f1��: �P �$Could not locate active partition
 �� ����t����f`�M r��� �����u�fa�f`&�w&�O&ff�� &��t� r��&�G<t<t<�u��fa� �P� �� r
&�>�U�t�X�� f`1۴���fa�f`�� f�>"f�6&��B�fa�              f`��rl���6�fa�������$?f��f��f9�wf���� r>��f��Î�f��f�f�� �������:6�v	0���s���f)�w�� �  �  �����Could not load iPXE
                                                                    U��c�Ӽ�0Ph� �PSU��t�G�� �<
u���][X�P� ���X�P���t�����X�f��� f����� ����� ��P$<
i/��X�fQg�fY�fQP1�g�XfY�fPfUhh��fh �� fh��  fh0	� j�fh�	� j�fj jf��f�ffnf�f
f�f��F����F!P�fV  �"��� � �и �؎������� ��$��"����fV��f&f]fX�fQS���Z�rf��fѻq�L�f��f���f��f���[fY��j@�d� ��-P-� P��d� X[��fVfWfU���f1�f1�f���� f]f_f^�f`�f���f��0  fQfWfVf1���f��fVf�� 	  f��f��f��   f��   �S��BfYf)�f��f^h�Ph� ��4h�Ph� ��0f��u��f��f�f�  f�  ���� f��f��f��  f��  ����� ��f_fPf��u*�����f��   f��  ���f��
f��   sf�   fXfWf�0� f��xN ���� f_gf�$$fW��f��  f��0  f)����f_�4�2Ph}�fWS�i���[f_�2�8�6fa�1��x��`�f���o��W�f���f����S�����
Installation failed - cannot continue
 f���f� 
 
��f1���g�E�ugf�egf�eg�g�Egf�E�fPfR���f��gf�T f��g�T gf9Esgf�E�ځ� ��gT 1��gf)Egf)E��g)T B�fZfX�fWQf��f�   g�G������f��Yf_���Q�����������Y�fWQRf��f�   ���� �� �0��g�_�]��Ј���0� Մ�t�f��ZYf_0��fSQfRf1���f��gf�Egf�]f)�xgf�]f��f�Ҁ���f��fZYf[�f1�gf9} t&g������g��[�  1ɀ�vgf�Ef��&g���[�g���y0Ҁ�r����fPfQfWf�߹ g�E gf���gf�_t gf�_��gf�_g�E
tgf�_$�g�E���gEf��f_fYfX�f�   �f��gf�D��gf�\�
gf�\���gf�EfVgf�Mgf�u f��gf�t7�f9�rf��gf�4&g�f^�fW���v�
f��  �J�g�]����r� ���î � �F�<r@f�ǃ���������f����)�g���  ��r��f����f	Ǳf��  f���&�f	�f_�6�� gf�UN   ��ugf�U�   ��u+g�E �	�*��gf�Uf   �u�t��gf�U~   �e��� f��  ������v����gf�U   �A��.�gf�U6   �1����~�f��f��gf�L�gf�f9�w(&g�$�<�u�&gf�f9�s&gf)^�f��f9�s�&gfN����f�f�����g�0ù f��sf�� �����f9�u�f��t��fPfSfQfRfUgf�f��fV���f^rsf���  f��fWf��f1�f��  gf�gf�}� f��  g�f_gf�} g�gf���f����gf�Egf�Mf�    ��s��,�fVgf�u ��f^gf�f���  f]fZfYf[fX��������    t��,T�i���-�|iP:�;U�0ZzX��`|@����U���9C=��FMfM�u�;�<�Ti��C7.-{ln�(+]ˎnii�
0��v/?�	8�ʀk�����;���U��}�V���k$?�CѮ�<���8���ۧS����i�d���9yJ�W�.�E�P��S�Z�q�v��&�X�SZ
����̐�~�>V��c���H���@���"�����������   3�X�Ww~����YU�g�$c�8���d[�u<g�%��r�������T\�|F��L�`���(��H����P2�"�f
c�-�_�\��>^?}j<��]��eb��u���ۀ'�A��[N<"�: �j��?X|=���xaO8q.��1?8R*g:�
e��b�j7d�s�*�3��*�Ρ�,��q
���LK�My�B���&��(�Һ˾	��\�?*C^��z(P���k#n$�i� �r�����w��I��#�����3Q��]qL,����f�j�;������㆗��Wp�[
�m;�X N�x����y�R�ￕe�E����@T]��F�,| ���@���%K0�ڶs���=<U^��-��%<ܮd
kM,�H������܈zr�ɧ�[�yu����S�C�)y�m��k�A��_��Y�G&�tf�k�3Q�e�Bi�u��_���M	~]�x%B�ٟ�r޿դ���u"
A�[�x{��tFEɹ���}�K	����h�������QI�@�40̒�F���`�:�,�FY1m�O�K�9�����y��x�"���!W���9�n�S�/���oX%,L�Hˊs�¸8�ݲ.p�x��6t���~O�^ù���m_��D��T<}�֮X�km� Ɍ-r��l��h�Oz��@x���/���^�o�V,ɖ�����2�3q�I*�>IH��#R;4��T���6�K+�v]�� s�O��{vՈ��r�;���J��s����	����G��m͋!)�T;�}�����)x����mZ�r�q� YK����u=�Q���Ϫ&f���%Hi��"�38WcH����=�t(sq��#�!4�!�Y�����,D��}�zz �G��_�r��M��?~A�G�\;�K=mL��XfM�01ʱ0���t���lZQ߀��w�����oA����{2�U�CĆ�Q	���S �2���x	���@��2�5L2�z���̓�_$W4+c��E�-3��O���Wzp=Hǌ��\YD ���h��5f���U��3Ƥ�1�%M�~�LUd��MȔ��w�}�tG��XQJ�s�#7��T�f�*�LP����f,	�li�Yx�UI�n�|�'VW1LT�� N��|g�����>�d�����'I�^��6��IqD>��Q���z����7�d���Z�aPJ�t�q�O��{܌8D�4�SN@�^��ϔ
l%=*?bj'm1�%�鶧o_AZ�{%6Fi��>�P�pB!��^D/�aHzY�o���e�UM����y�I�Т�uz�������5;q��`c"য়�ӧ�v�����p�[���;����O�>��>Z���̠��w|�,����8V�����=�T3�T��X�:6ŋc��1r�ܟ'��5<��h��?�B!k����97�x�Pm������ap�����&������Dsr����삺���4C8�E��h�-U�]��A`nHm|���s/r�V{B���n;��z���r�'��������J    Hvπ�㖞�zq����v���vu��M��{�qz.B��ʺm^-M'�X�M��=��t���K�F���MS� |Һ���  H#�%.�D��׃��D�
���dl5{�&�ܕ��cN�Y���Ռu�+�3�6���Ғ�[S�?H.���4��y_��ʇP�|���cf�8�P�����\ ��iX7N'�l��2D��f�
�N�g�h�7d�@r�
������]ƛ��H���M�m���r�Yqb^}�i���W�z�_�3
D��2y��\��H�	��7��#�㊑��#`~���e?�$VK��k���йIY���VҊ�q���� ���v�rJGo&��rb���A�qYRnm�� 7�Tsdx�)+�~�SI�^�u�	�+�纖3�c�2}Yw�U�}S�T���Y��TW���R�9���0!5�{_x1!�}iy9��&��
a۱�����D�AG��_�v樔I�_�:�3�鑧(�=g�"��uf���fC����Qa�+*����{óBkq�V؝��+�2$�*]{�����	a��6˭1ڿ���I�
0n�m��(�����u�o+��#Y�Q�_u�-��g<>�!��垉8ы�|io��d�ڜ۪@mN���uz3z#pA� �61�"]NԆ���DniT�p� ^����HŜƷ��X�Pٮ�h��%	0�n����p�E~$.'*_�&��6�}���v���������k"���hɷ8V*�)I�pU5+7�-����(Զ�P�,%���Q�>r�r��{=�LE��\�A;vY�0�JaQ��S��$�4�®"�t7�_=m(���2_��n9hz�0+Dyuܪ0΄¿X�r�L�D���^�x� DB�':ަu��`�p�6h�<#0=Y�e{���8FE�ɵ�O�Ex��][��_.�3�����Xgc������9^�j�������B�c�H^/�qg6�t	,a��¯oxs'ꔊ��W�pT���p�H	+��y)��M��exo�������t��h�t�����c�<V�	X�<L.����'d]"�C�3��,�ZӏR=�P@����鯲'ɂ�Oo��УfeǵK�2Ĩ�����M��nX�C��f�� 4����6ʳ���L��A��A_dzu�{���__�ލ�u�TϽ���L�ɣ�q�e���ca������m�}�f#�d�.^��H#.⡔🡂cV��f�"���8������*�j/`J�پ}�p!�T��t T7�yi�E�'�L���WA�e�n8��'��_4Q�
��� 3`�� l���&�|�]WȰ2��c�����q��Mhn ��΢�F]�V �h��LV Y�qە��W��A�a=��<z��xmg��f$B�$L�s�a�ڳ����%^�Z�;�7��H�M��bKxP���!��}��E�Zc��3�Vܮ�.�$�q��L\�I�&!���f��n�WYF�K<�3R��l�g�������`����`��Kt)�<
��$���?�M&�+�p �����J�W��8����l�ꄺ`���d�t��a�t��ۨ����lU�*�5*����is���?UE{�;B�چ�=�!W>�e�8ǘ�4��kZ�D�ܤ�[�I�\��}.�V��wis�்�l���$��MZ�ڲry)`�ԁ���nc�̈́}\���<����9�?��c�5��'�!Bw@R�}�fN]��Fb��E���7戥�S��F���\[�Yxl��>���rո�ᕤ�;�gN 5����{���^��.+-p��k�����>g��}Z�@L~/��Χ��3���� �"R������K�U��E^"�&;��rx���a-g-c��&�iuv��:��"^}ڗ�ݝ3��hk�CD3[����{Ēx�z���&
�=����,�Ko� w��u�3�p%�w��۾�^ۜ7c�b\������爫Eui����a�"*K$3�j�Q��#@fGîa����\����K2��m����� �������Ø�6ȓ�|k�Ҽ$=��'>�{�(�F�VM�!��W�Qa���[�z�-�1 � ��������a�q�)��8��^�eo����a�{��r�W�^o���"`�9Y�uJʜ��I;�W�lV�������,������1D5k)^9�&����#��KB,$�_� �A�S\�~����e�)��p�@ z�$�K�@�IeߗpD�Af���#pB=9�g�A�fr#ѯū*�,4��K��wVV�B��#\X:`��$7���}+>���~E96�ьO���Mm[6�<�J��*v>C��=�*0K�7#�?5w4�.P�t�s��P=����Ȥ͘�����A���
E��U�2�(���51I��8��,2��0��D�f8����^H�b�p\���[Y��?V�qnYi2i�Y�6��FM_��?oP*��D�{�Y'��ٴT��&J���b��~��$Me���'�ǝ��K1�0HP��I��Q�υقWx.��|��#�t�r�{�c��X��X�N1��K���0�f��ʧ�_�^�c�k.�%5�3%�9ZT�:���J�ԙ%��$�˿��WrR3eDc�悄��y��3Ɍ'�kno��Q1����,�"��0y�����Y|ng�z��j�T����/�яxAѵ�ҋ��!h��U:S|8	S��G]+����=��̒��z"�i�R?�&�Dn�l��T��t2s��2��w������g�����8��z4��������.�Ï*8�>�fz��1c�S��d�Q��vd%C��v��E�f팫����^��U���9�7�_p�C�j��P6P�u�2��N��8�괓�����WqR�!����"�U�1KV:����X��\��@��-��9FS��_���(�DD���ў�ř�t-��Ծ�s���TE�&�+�?kC(<쵂��T9!T[�A��:���l��{`j�뒛��h�.�$�#�?y����
u���lJqI�B�d"�X>�6�"�dI��qk�P��P.�К΍G�jy�W� k�:8%��;|Ǝ�&��4�F��{��Ƅȟmʃ^fE��瀖�|m�����0���ZV�=�f��iv�<zbQfnf�G�_�X����P��U��*��څ�'��H��I6gY���v����֮����vl�w,���A)�ݢ��*��aubϝ��������\ό��q�u@�5"��N��4f �8Yn�.(f^}��D�M������z{-�0��e����u$�t��{�]����k��_�z��Qx�>3��KJ°ϑ+H�� _$�Ӱlo�b��S�=Kw�u\[ܚ�O���g�8��HM�G��f���8���8�ݕܵl�4�.?�$�SFwj�>��7]{�b�Z{�����L�\[�z�#�p��H�vi�\������e$E?D򪾭[�e��H��Һ9�JMr~Σ��/3����O@.�Bֱ9�
iݠ|S�j-H��D���X��'�C}�1���� ���Tk%�:)H��F��b �x�ۢ;q,�k;d����n���!�J� ���]���0�m�B�֌�����3�?a�0�>3���j��Po���QX���U{wN�X��V
LXT�v��#���j+�IqnGeX�m�,-��˴�C�;wECxdp.|)7R�}�I�%��)`_�+���"l9Æ�E���˧&�y4lh�JyR�h�%�_θ�T�UO�E؂��[��,��g�L�'����KL�E\3��z��y�#a^��8�k�rJ�$��w��OuGK)�9}���A�W[�OJ%�GW˺߇�L��T���o��*����]�/2��q��]p�}�?]_t|(��RGO ����V�^�2����h����C�J�6F� ~a�ȍY�~)��=����AҮS8���"���B,홳x5X&��45�=Ǒ����3��E�_�3����`
B��H+�{PN�r��{2�O��/���敇���^�m�t�,�G�=bܝD�Mim���[٬����:���B��0#�y��E#_��w��S<`�K��9����,M0��Qmʫx$�*J�#֌}��KHl��X��ڀ?���*఺��]	�2�N�׃d����hG��LZ�!��	%٪0��TO�Y|"�я"}1���8P�F����������0����:#����!h�o2�~Ap��'u���]^���mθ̷*��f yGN�ֽJs�YRX՟6�-�.l�u�4ڹ��!��3�ȍ�A�S�<y8-���?��:b�xW�� � ���d4�Qn�)�!�۶s��3��Z�4O%�S^�e>�>?�rs$yZ��Ȯ<jp5����2���@�:�#ѴHǆF1V �qH��&�@��G�� 8c�L�ٟr�܄0�j<N�f�RMŲ��G�?�{𐔳������34cX�2ǭ�=j��g�u)ewr�t��E�2A���7(�i��s�m%h����������4�9�˒�Q@��E�>�$���J)�<pw����� 'W+�,��"g)�z��m���C���������Ș�T��	I�T�&��ta�S����u/�Zw�P������V��bn�:n[	42�׍qP2��6n��H�}�E�gȷ� �W��
����v�]��G���"t�qxg�y�w����~�|�7.�q+�l+6�H�',�ڥ�5 �A�/�.��{@�;v~�q�Ot�@���5���Pێ &�$�S��n$�n�6!�a�a��rn�i�=ѿ^[�c-�w�-;.:�E�q�>8�f3,�*3ջ!O���KI\�g���e�O4�
%SR���r-��"��S�� :�=�@�|�;�c��ESg'!��J���o�]��y��Yc�\�)�������Q��ڲ��G.�t/��;��س�+#T��R�P�?���!�~x��X���2�­O1�K��8j��d�R�y�z��7�!�|�]9$�=U���M�k��Hg�+�P��T/�Ζ��>��0��C�����5^�>b�ӻ]@�9�ܰU�h/�[�|*��e�?X'ȝU۲�|k�b9�?@>n���+z�P�t_�z�������X�$0�.ߔe���tmI���Hf�;�ھ�ߠ�����c-���hoz���THC��x&��	�R�=�8�ɹ=o����)Z����S��9��?P!�#�=o�>PH�BB�_r6�y2%D4L�fhs��[\k��[\y�4���D�A��k�.�ً�G"e�p/xC-���v ����=���{�N[��Y�[�$E@����/��9�=9�J [/�s:��\b�3iY�YE�MȢK�ɗj�>��J}WTw�L�O�t�iu�%�:,#��Xƈ,}[�ݕ��8���KM-��1i�e��� �����L�y�Fq�Y^9��(o���<�>U�F%8w�Bk?��"��u=�o���Swq�V�-K�]�k���eD���Y���8�
��qԈ���X��Q��p6dì2��z���[��ʩ�S�����4��U�$C��8;�'��1����V�D��z��p�䚍x]I�5��9��c��ȻpywD�S��۽G;�x��6�p#a�62o���G�σ�ӡ��m�Z���lGi��*���I����u��6�@#�����r�H�MYP���W�AK\z�S���^޵���J>�ݣ0������n�Nv�]�H��=k+q�	�}O03�o�����g�:5��S�[���ӕ|O���CO�P����σ�5o*�����
�����F��Q祈BD��H �cn����L�}���5P�媻�n��78*����m�B-�J5���=ǸL���'8o�$���{�����Zm������kٜeCA�{^��K�8��P����0�.`(Z����*U�i�_�I���R�R?�	B�S�cI�a2��g<;�f�#�j<��܁���I��Қc܏DN0�竮�u�$<E��g#�����Z���б�KǸ��5����FX:?/�%���N����
�!ɕ���Ž��_���◗G��?1`�A��Hi�fZkkW?b�g�QI\�F����X1����g��ם2Vb�>}�/Kb�$/+�u@��GG��:��Nm�o6Rm�Te�����R����h��2.�V��+4i�/9� ,>��ǴH3�r~*��ۄQa�Rņ�˙&���W�1< >K�F_gh}[�dB��گ���ᮥ�;���YF����wq�Aį�����3��;�緿�G�:��f��v9�J��xW�#u6��i궉d9��%Xc��S�'[j���~����\��;�|�u�IL�'7��O�����Q���&eNjҨv�c�!�JL���}�?c�y�/YysoXZ(��lU�}-�
V�]R+�$ڸy��;_v�j�_:#�yw��]_t}������,�{�V���h����G�����8�e)����$��;�@M�Qz�+FO"�n,��X#V?�S�cq�+�zC�(E�C"�Ԅ��ǀ� s��LIv��uB"�PC���o��t���NB�MS�	�=��+z�*8��S�?B�Z�\�N�%��o��YB���{~;(�q��&�4 Y�׾E0,bտ��X�T6kI��%l��	J�|��꾯��6���c{�w
�{t9X�x������Gaö��ok�BC�����F��±4���<��"��{����0�dz��oJ�櫝�*��k��Hw��R��' gf�1iw�5�@"��h@`�8����io*��l��^G���s��dX��Yl��O>�/��H~Mg�\˟^{W1�5dz��
������/g�t��}k�n��G�m�]Jf�Y$!D�i���IE��`*b=Z9��/�\�o�K MVл���5{h7OI�U�㒆bI��p�����u�^�`�ZhU�r��f|�ާB��=s����FDk[�ozf��V 4]����|s��Al��,6t	SDvԪ�mX��̙N��q��c��_S�N�wˈh�z��X'��f�����Ki�+FC��C��
]{�����n�ۨ,�8�qc���gI=E��!�߂�c;�9��A[�V����:��[h����1��;�0�ȏ�U[$��7�>��/�h�GFCSo�oV���b@�US���_#�Ҙ\�ta�y��L؞���o>�*~�}����i�e0��2�b��B;�/DdQ�Dj4���_ꧥ]�(��Z2A*�wT�kbI���"c��S@9(�(���n�,_�[�H�T��k�;���m�D��i9�a��{8�p,U���������)�ȕ�r`C�ud�4j��|P*{�������S��8Kt�m4S	R��~<(���as|ܨ����񜍀�bF���2��ƹ���Z����r���;���ɺ0>a������L!��-L�2p��N���x�����j%��(��ק�-	���q?�c�w�"#�ƴOO1G-DgW}а�>���Q�!7���v�u2w8:�Օ������Y߾��y`��7�FF�3��� ��d0?!v�,f�Qj����ܡH
��g/&z�x�a/�	�F�F|���{�(�S E�CǶ�i����M�A�,�^cOY=���f�V��'M��af�c;�PO��B;G�"B�ڃ{�-n����U�p0
W���a(�*ͅc�\�p���y�b���DDk�v����jL^�覈x�&~`��Z���af�1��������Y�ҕvJڎ��b��u�c�-�I��E��4*XX�����Mq���(o��b8M�%p��bQ�c�%�
��כ/��^VӒ��}��(�J��iK�	:uL-�
JUa���Eoi�M����P���|�I��paձ������^r�=��0!D��Y����=��ۤ�xdy�TUf�H&׳�5�"Kx:2�K姲�K@hx8�N��bOC�-�}�r��F5n�K�ط<���o�1���H���R�V����oA[�G�22�����@�;����A�Z]��H6q�'_��ͭS�0	t<ä�C�:y;��{2hQ�gF~A�$����Gq�Ğ@g.��B��p�z��=�����]��֊��E~pl�o���=_g��.S�g3�z�ۿ9+u= {�ePͮ����7�UR뭉2+% 8@N�l��A�&�·u���+���f1R:OeP�9���{��
������W���������A/�B�+b=�2�h�q��l��� K�{'|8�M���XG�<�	��
�s�S{%�=�z-bT�7J�eŔĕ��,#ivb,r��9��ʠq��p�~����Q5eX�x?�ע�%��:m(���r�����?���_�X����lgäp��(-/�r����������L��e&�}�[!�bi��G>�Ƿ�[ڻ�`�����t#>�#!����ᓍ�	��r��,���`!��v�t�A=,12ʸ�C����h��9;�<m�0��m ]j��u���qw�%p����y����6F�����*p��:<ZI)��+Н�>ӍR���U]��q���I� z�z?����љ�F��U�r���Z�.*Jc0-���;agn��_i�\�?���hn~�}Oʔ-��fŠ������w*&R�M����5,�+��m;qm@ӿ_�N�8�����?����Mә�ґ3w>���Y&7��G��G�{���i���2��w�_g/q�^�@�щ������P��q���C�+��R6SB2}!v���I:��io�2^����ͮy�_\�&BX�- �ˋ��T&X���^r��*�Y_B���M�d��~���8��c�e�~��L;�	W(�$�?���/}e�dĉJ���U~��<�����W�Ny�m��X��j��`�_�uBOSu�	��_B�̞1���~�z���-����Qqrބ���3qqk"���j�T ���m��8g���V=�(V��D��ё��A�gtǵ�^�FL*�^�GV�-R|J Mo �4��/#e�8����2�k�u���O�Ex�6����̓�ҊZ�������k��&�p<�ٖ�(g/�T.,�*�o�9Ȣ�鳘R���"�t| �+ϡ��Z9-J�c��]lm~���!��|��|�1g������J-q��1�rp���z�����s:-��C��gm����5<��$^��F�Q�u�
)�{mRV'#�%=��%=�m�O��v�X}p풣D���>�z���C��V؍� ||�S��⏤��#�r"����ϰ�o��Z��;��baW����*��2�!LCc�D�zh�$k�2&��/D�����L}ar��w>E�,�Dt�d��A�D�|:�[4Q���Y�^\��'P�)t���!��G���'��Wu���~؜)ECǥQ�S����k����#�y�&�(�t�����>?�2��vm�&y�K��n���;@���.(������|8.,Y�������Y'9^����p�w--C�@�bۃ�/"�c�	���S���m���"&�K��ל����l,〃[u/�s?��6)���!����0�5�M��o.�n��ġ��'�G����>�^��EPkI�?&�=�0�)�b�ǁ:LD����7r����H�Of�����:����
m�𥑋�$<-�O�� l0�\t��v9YD���Fw,5���(�����l�:m���3�j�A����b��LeZ��ǰ�M����0l�>rKX�$����r�\Bċ��=qƐ,�\l�pt�$D���O���l��YQ8���S��%7��p@ႍ���a�:���Hܫƴ�ɉ83ѐ<8�Pu?�mGD��k����0w�O6fN�!�'���@�v�d��cϼ4��ngV�� pZ�z��x��nF���9�W�����ed�R���LV�mX���r���6V���`3�@��+�Naky��q�X7�����"�e��^Mb����I&�a�����1�\-���VTw���B�T4R�튡�ۻ�X����=�h��Z������k���W�7^��r�*�B�{����Ϋ���0��:����ݡlP���h�!�6�O ^1a}Hr2�x��'��3�.�o�.�aX	K�t⅝@
�)�Y� �ġ/��Β��oܡyi���o?�o|�߽��;���ńH�5� 7��5���6�����s�����q��tWu�ecY����S�80?�i�H�����m���i�XNZ��W�#�ݼ�
�<_.�`s�r�Q(r��d*c�@4#W�/��ɑ�Q��g�s�U�U��]5�TTJ��&����S˥�#t�j����;�e��>��[r1P?�Kr��*�2���Ʌ���|���0ĽT���Ci�6|s��"�*n���_b��;��"�P](���['dw֯�1�%ͤ��Oc�H����f�Dpp���'l�;�e�2������6�l��EX��2r�y��*�'՟ىO�+8ML%���Zj��U�hy��zˊޛ�W��(���5f�oiMG#\���d �\9�sT1�-�U���1{ذ\�q`�^��v�G�@"��5��4�b��Z�(��md֋�����'��X(<��)�J,i��_��K�����O�c�7X�q
��$G)>E^����e���92�M:R��P�� ^M��Ohs���6hJ�~3 x�#k��f'�L��2��T�Z�=�)C��/L��Ｔ�`��r��֜Z�ݬ�۴��H#���ї�>�����D��f"	�)�@A��7܋ʞH���ݰ��!R��)b��C��;z��YU�sd�Fa�ˁ������vz��t�:�KM��W�u��P:���
��Y�z�!�+�(���D��'1Ҙy�"���W��[H+U�����)c�pY!4@+.ps0��Os[l�շ<;��wF��a_�Bo�3S�|D����I�R�A`����4�� n���d���ۻ�n\wA���/��~<�h؇9g
����� ���~�����A3$�bS	rẍ́ة��F�����w�ΨhG[r�v�~L���t��)�����0>���}�m,}�:�~Do��� �kg@�}��k������������5�kV�q�'�7i��[� |���3��{����a�x�)�7���� <CvJt �M���@y�P�t�~��F�O"m����{i�����+{��)�}���� ��P�������6
ث������\�Z��;��(�?�x1\�+
�gcb�5���1�3��[X�d�8��X5ɰ���lV�	�6#�l���@��ͩo!���F���Q�S�R�Z�?��C��0D��psb�X_��Y�T����Iq�\�ɇ=��T(�Z04{�<������%�~9�կ��3��a�[�=x��:5���ǯ�����ǮR�.tO���2��.}�.0�}U����x�{�,����E�q�\�Mi��h�U{��"�U%b'\�;�x#�fӜ��x���e�M^�]��"b��X�׍�ex���@��遟δ}�k�����T38���Z#C%eB�;	3�S��9�1�����O I�4���/�+M��e[�L�c�,��(
��%��^""9i6+x`JR�����_�I:�vB/���@8n��Cப�j�VA��U�c�Ӗt�.��
��#;T���Vt��."����(���>y,H��Q�W�Jn�ET����ܲB�:�n��Ye�U���&]=��#\b��Nٞ��[<����	��'����|��@4���D�A�]e�]zz吪^��X����B?��6����H���gb���s�-���4�w���ϓ��Œ�Y..�^f$�&O��ܽ	����lu��W�L�ϞùR�di�Ym[��}�OFN��,���)�A��V-%)-�)�1�/"d4����R��(��}V�?��iZ��v�;������Φ��N��!m��e+��gN	0Ub�n ���O�!���[�qh�V}��p�5T�~ܻIL]�c�9a�[����B����͠]"p3�lh��Ҟ���;�i��^�,x��#;$�����s��q;���簄B�� 5���騀7�5�^��B��K�k��]dq�`�V΢��j`̊d�wU(�Nf�F��� �kW�LS��g��Hd8$���_�����[���̙�F!Ht��Vj���92�>FF�ڇ�~�� �_P])�A�(�!�I��2; T���mH�b
���27����H�R�LM�|�h�*�^���.�&6.��o���,�A�L���^��y,�qT��VL�����Թ�D���p��2
lGQ٤$����Y�w_�����(��2_S0&,�<֔�d��Dj��d�wz��5�:����:�w�s�cà�[ӥ���ۭ�0�8{%�抧Ѱj��i�RH�?��u
pRC���.*�^��Z��	
	T�b�۶��~@R��8
Mީ8+�Y�mֱ$���5���%X�V�e�v?�L���^�)�S�������|���*�B��r���w��&}R���-Cm\	��2���iC��H���m2��=��% Jr���jo_�G�<:�pw���E[�l=$�A�ؾ8z�b!?���͢F����6�.'�M+�σ��9y��=��&�U�~j��xG�h�**������&D�J�dW��9���/�B~]P+8�>�o��x<�kI���u�3��#�$�P~�2u��۹��M���l�rTl	��˸E��
��N�@$�(��~V�^��X��XAٲ �)|�P~>��������ll���K-,3�?�d�~���G{���UGf�Z��p�����@8l�����w�޽b�T6��;���s��7�G4^�\+	}��(��<��gX���zY��ۈ}���:�E�m���P�3�����O(����$��Q|,�Z
�AI�v�~�f�g�j}b9�� �K�"��e[��*V��a�����(��3W�	�y��V��`?�ՓTL�G������+D��e�?x*2��
9�m�Y����O�Z�f0��S���5Dq�ӟ��F�Kx��`r�|עd���P�A}4-'"��C�}/�&�l6�k*�AX��-���Y�*�$W�.�����l���(oq�~mD�� ������uٮ֝j<݌#����$�|�~���������'�$ ��ul���N|��)݊�jΎ��:�?{�WЊ�m���'8��|�v�е��	L��w��^q��J����i������fwҔ�6�Y9>	�R�yu�P�1p������uB&�1x�:�ĉ-�)\��6:A!�ߏR(�.Y�]ci%<Z�:������0f�]��+IZ��@bV�&�k@{h��\KI���yجR�3(80j�W�1�i��Ȉ�ƌU��$����vE�� ,��}3O!�!:P����'y�Id�L�!CǍj�:�j���OSA�J�,��ņD�ׁ�5	�,-���C���]��ML��.6����wB�.����NG �A �x�*Qj"?M@4��2�E8���.&�=�*c�K�9u֔@̮��ka�������G
'\��j6_��M��˵xB�}��R�1�Su��B�Ӌ����Ş6�`F8z�Ǜ�����2�Q�<��,8�>w�T/���5��Ak~(=c�+m����FY(2��"�(Ϟ����/�a=c�ލĴ��{ʨ�|�i��z>y�M���j�3=TGa�����$�.� 4�<��8�_Z��9N�u��AT�)��Y��h�Fɀ�P�PmE�w,�%�U���]�|��:Sq�hx6,#�U�yw��O{��
.]�g^Q-Z�q�{�q+�p�}�Z�y�M
T���-��H�C}����ۀ�J�d�!�5rJ?DV35�C`R��E�Yg��^�g\�dI�AF���ra=z4l�̛ʹ��k��6�'��C��M0�Ug'��"���l�֭jj]SE_�-�ee�_� �&�A�ceL56�!��@L�
c׻�ʤxi������њF�N���"I������ɖ�l���a�δ�S���YbO54����w�a#7�$y&%�&\�nK?����¼�����в��y)���j ^BR�"K� D�F<0����RE��L~?+��޸?�1��� ���I�o8���	Җ�F���!	9��W]Z�"I���5�,0l��˨P�Ԓ1�o��"���e��S�J��9��E�WQ��ʸJ��y*�+Ke;Y+殺��%X�Z1W�ӄ����E�s��A2GU@F��P�z5�t566v�����B���0���MAt�N�k�Y���g�ތ?���Q��Z�:\����XR��`�a�d@a�A����*�'p�H1aP�W�K'�'!���1{3v<"����i��R"��;[��)����:�$I��v��1��~��Pԧ���Ey�>&[��X���ǆ�z�2X^��\�F���X\�R3��q�\mVt��	�t��9,�.�|���`���[����k�E���R:���(١C�L"���n��<_�������K�|��T\��V��B f��C�$C!v:��|e��	�s+/�0���J7[���"#�?OSc��{.3��������]1�k9�50ܛ^��7ڟ@��R��a���X�6�#N����m�;�WP����I2�X�O�n�>;>�F�/����b���\�b�@��~�l�a���,4r�Z�a�&��[��0A0ƍA�f�r�Ys2�\b�9��{��`<v�OX-�����9��)\fy)����[������V@{M%Ι�ۍ���4a!Y�Tq���Y����p����d��}��h���0�`��{J�a�ȋ�.V��v}��l��
`V�e���4h�}��bI���	���i����""�N���(ԯ�(^���xPy���_��U����:�p��y̅�h8;$ittX�w��T��p� ��DA�A��qR�˚j�Qc�1�ɯ���,9y�P�>J�r�GLaDQ�U2�ٞR�m�?1���j�ǆ�@?�S�*;�[eE����h+\Ys$	��R=��>�}V@������^��
yB�+~E���tΎ �֩k���%;�8ϼ1ɶZǒ�i�ZdB:6�k;�u�W�5@W�֢x�����@)�ι�M�r�Cl������J��y�V����U�U+��R�����?ے��@@��n�a��u�W�
���8�u)X{�T�+�ݠ���C���;�A؟����{@�27�-�ݴ9��D�x�[��/y�u����?�F2(`ѷ� )�z��A^�i'Ap�3@�N��ܕ��Q+E�+j̢�1�cW�x�ɦpHV����<��z��x΅�]�/�z_�l��x�X��0�+a���PW9�}A�q�-���k����� ����$�s�!�N�^��0��dX�x�-�Ɠ�c�y�U@ታM�5a(���ÿ�j��6YG�W�bP���V�*o��KY��H]�bܑ�\Y
Fu�/R�^3c=��A��/�h#���O�f���� �U�/�R�K��?%�L�w�������~�S�~�A-.��נj�*�n�#8؏�5��#�9Z��R�F ���tz~uJ��-'?M��d��Ħ9Н��l�j���X���Q�Z!J
2
�.-��0Qk���xF�l�\h�R��жL~������"��j����@fW��L��2�����a(8>H������ہ����N��d�7�zJj6J\N��r�GI?vq�|��߬�3 N�bR�1E�١^-
����.������W��W�P0�2�\Aј���Fm�a��*�b�ޞ(%`˗'�S(O)H��nt�e�X*�*�cr�1��b&�0"T�L	��R���sx̀#rXuW����'��N�P@��$�?���`evqp$�FF� b��p��3��~VG7LWK0;gm�Lx}~x-
�,�o�`�8m��K�q��8�-���k�n3ZUP�h^&���=�OL�%@yqʶJ���$R�>%D�wpU�9۪����="PS�o�oz��X����@~j����=4o�g���6���6̞�RM"��4*��G!������ZQ�n(�j3���!I�4��{,��<?�o��MNy)���B�|_�nVyxj����i��������`̌F�����]���N��_&���lȊ�M^F�Κ�|	�!�>�i��MWȚ���r�a�ȅٚ(����Fk�S۫JT�!!��Z�)�H���#����~#a�ݙ�&�=�;KG����E����x3��I�����UTg\p��O�,�9�W�%�mۑ��͔�=��d��m"A��(��V���R��#��S���wb
�篶�1S���:�Ǚ-%�5w�,�WB���heG���g�AZCx$ӈ��OK��g�>d0��]�����Csk[�F3 �rw�l�*�X?�>��$�5|[�@�:����A�_3�:d'�����i��`	W�V��!��zk!qw�H���]Y[.�[g.�b�*a���M9�x�c��8�T:|ʯAX�ш��jBLc�V?`*˪_!��wy��C<5z�t����V�j�<�b����j0�L��=ฉ$N�B)z�tV"0�����,����E@*���f��k�ViQ8U�06v���׽AH��y�ȧH�Cn�/�'n
{�-IB����,{b^P��p��D��'?,�"��e������H� 8?b�ս=��������3M,Iه���M	�O�m�b����ԥ}c���&]v�ON_��;���~'r�N;����';{3=�x-��'`���p{<���䖩�c������4Y�V�u=8M���؁5b�����f�WmX�q#v�+��l�6�s#�뗯����	���8U%:,�����<!&�a�(����)��+)�5�9��k鍿\��(ď�)�/�G��"�`��h�@���%k$�M�`tgٚ7�+��#Ϙ|�t=�{�>�e�N�8��S@�B"Eౢ�p��*���������TY`uǞޱ���q�g��wnI�E3[ت|k~�I�2�d��	�W��y0#��4%!�Κ3�]��Sd�����v��/h^�vTaЏ���h��^ש���wY����S�X��1"�N�U��M4)_��\�D��u�B0\��]�����9�:����L˲� �l��j�iĮ��Bt��Yjb�S�i�\�h'z��Z�"hǗ�e��������v\��{50�TY��-`H�Mc�鈦"s.�JV�)������˯��UVOA�p��%e��D��x�q8���!��B��h2|���K�Ⱥ!C����H�-�-oť���W�yp5�;@�/�h[lX1�l
�b�V{"�����b�ԩ��6�	J*g�y@�CB��0UYb��J��4���ۤ���y`��#q��A�.�����omH͙e�����|:2+���ɥ��:��Nu�Q4r���xcTx��V�f��,��\��7�ALxJ2-�P��Q��T�lP8-�7X�=8A��C���m{rk>+�N,WYXJ�2Z3c՘/Σ�Ʊ7�/롢t`'�������JxyX8�G�Erm������(�(�j��(���`TyOG���
���`w�g�g�pj�����G����� �w@ K���� ɸ�!v�ݩ4h��.�@�j�뛝h�g���i�P�����ʘ����1d2Gs�a�A�ׂӽ��b�mV��w�&�D,��g��Tҍ��W.�80«��l�<�8k\�@!�']F�qYF鄁
�b�eK������|LR��W	���Z�?�s�㓳 �k��>�ʃd�!h��RMw"��K�U8g{��f�5�|��82��s�i��6J%��+Y��d�<a��U���4�Ag�5y��b"���띹�f���h9��m�y'�}0��l�6���id�'E,�tk`�nlG�
=�+�E�~� 9��p�N�a��;^�_);	E�1�u[Z]��G�*l�D7ⴚ�^h�u�=L�%4�u���r�E���nm�[E��U��'��#Iѭ���X�PC�E��5�Gx�h1�@d��y���P+���Z12?�y/�����_���ƞ�Qcُ�m�}��{�_$#B��K���e>>���X+�3ēf��uRX�N�WM�&���6��k�[��1��|B3��gc�o�3"�N;,���j�3�+�{�T�2�U��=#��w�����E�F �k�$	�:Ae����T&�`4������6�mMj�7�������&[v��+�AZ�&߽u_>9Ԫ�SbB>5�Q����~M啑�<�>�`-��|E���r{߱�����qŌDcmK��Fe�����n
G��f�S�Z�2��&>���S�1Bat��P�Hl�����V�W�y
�k��?�{��w��)��e\���*~)T��LgZ�3H㲀�`�3�T˒�
�;B}RA�UNe!����\��~���� �ph�L	�H�^ŋv�	I6�A|.N�6B8��ɤM�l��r�^\��ޜr=�M���Tt$����665����*�{I@���Fh�E+x&�[���8)�,8��+�BbVOJ���)���Bp�oȇ>�8�����V�'�Ȧ�5;��1&PcH���ʡ&��_��4-����*��k��=]ɀ=	�]'�K`HQ
�@q�?�ǖ	;�Zv���}��Nʎ�@�(��R���,��$=۝�T��(���Y}@���=�?(�I�8�.�\b(�/F
{W�z\Y����W�E�F�"�Y��3�=��QcZ��ʰ���Mhng��0DZ�\dt�d��m��eFYb����b��}f��э ��!5h�)-Y��s 	��U:��9�W�0f|	��kXR���,�P��魍 ��b��|0��C-��BG�J^�	˺�_�kRe;����5;��bW�$�lf��3-�!��6o�)!��ې�ڮ���?��=�s�{���؏7��(8��R�8�ŷ)�\�f��G�@0�cʬ��H�;Y��P�J�{���D��X�Ɵ��F=*�=���؎�V�җRaWX�� {����Z,^�b)F�C�g#�Մ§�r��I�{;RL��AY`�G�WM���� ���1�a����3m�O-Q��ޜ�w��`��'���/!���w&�Z��������fF4Ȯ��3�����!-!��g���i�/��u2dA,e�s�t��\�֪�a�󁫉' ��#�,]f�~�$.g�!3h��Tu�>��ا�ӌAQ�=/������.�=EeE�ϑ�Hl���s���hb׾�& �����A{,~_�k]E�@B�V{�Sl�>'�+3kuk��i�J� �������V|+�ܨ���n�Ii������8@p&�zm��?s��@���QGf�+�nǞj���Jl������Z�2_�,�r[Ĉ�eޡ���!?��r�D��7$��)3�H,����?+p�����z�H|��P]�a���w<�X�4���I�;����'�^p
R�Fe�m2g!6*���)S���6���@V��;�t���cS����F|�i�l�W�lI
S��V�+�<�d}!�63oG�M�\�~���]ao2@k�'�7˘U"�Oq�1�p&��:KyF�����f��
J%ȶ�et��I�۸
�0W�'h_�_3�7�{�}�w�ͦJ �79'7)7��,<Ą��Jg0���>�CS�P��^�c�Nϲ!��eZ�|���¸N|�W& u�t�k��;�u����i�t{hD�a����fi�$EO�	t��3U�c�h21t�%�C�w���d|f��$��1�O��J�w6g��WXxѪ%���]�lY�x�AΖ_͟0���盕~d���R�J�&<�Y�z�.`�3w��g��H:�e����\ 2d� =��H�H�l˽�������\����2d�x���\��8 6`�?��D�����6�nՋ�#u_%~�./4oHͧ��c��H Y��{��!)
f�(�����͒F`�\[�8z%ۘ�7�tٹ� ���>f�ڟ�
��O�<8š�M�:�E�gB��g�
u���	�O���,�5U�moq���,�~Wc�שׄl����t�er�"�"7��`�·*�t����
n��^�nd��$Rm��F(��Z��懧���u�ׁ
"&�� ��8�I"���Dp���k�+��e0�X�8~�.ڮ�ɂ0K�0�l-n�|��2-?x��/PtD9kc�?�d��^���5k�+�o�#SԆ��f��f�5X�\=Ȕ��)S�O.���rmdu�T-�z���}E��<SP{e�H�qkA�'>����8��[��0N7�7]���ͺ-�������I䅯ܜh�w��k{M���E��:��i(��xSԌ���g�aH:��b��ѣێÜ��^�C��<AP���'��[3��|h��{��X=;�2'M�c�o ��.��c?<�[�gb;n�t �-��+�d{@�j@圉Ls����ImM'O���~pT�e�z{%H�}��j%�>��W ���Uǁs���]���؞����w_���������G�MW�"�8S�A}En�h��Ȱ�z�� �ʂV˖������a���l��^���1Q���Ӝ����U�-�_#Ӎbn��E�UO4��>���b�^K���!s�
�M(�o�k�Q[��'�$2��ht�!O5"I?�Nއ^�R��X5bWq��'���ϼu�A��Y���ïil-��������U������Nq��̡|�X=����z][�<Y� ��;v��yDZ�@��z�48�)���3EK0���43� �� �Y�,�N�?����=���#3�T��"�"����!��]a���G�W��[+�&.�*�4Vk#'1Ns��P�=�-�8|72yx?h���J��LC��e�#h3*	1溘�P]8��5i�Q�i:��e�/(��'�z�n(4y�d����;�7%�h¯��7��,h�3(��:���H�9)R��(���pA��揊��~�oz?�)�?N�q}�`#��M��(h�����)`c/(+-�,J(� .��v���$��#O�>�kG���{�uau!������ЩN��;���$�q�y�K��R$6ʷI�N�ؽ�l��Җ&ȶY$�D?ؑ�f���X���AƓ�n�m���FyvYa4)tJ=G9��Md��;L�L����2$��޲w�<.��L���|�;�Ø�$�I��>�R$1���W��	��:��� ��L4D�y�����j�Hl�۫�}�o�3�6`b(Di����	V�$Q
@>�J��������U��,wW^W^�W�gg�g�ڝ
���(��\Aj��C��g���d�lt���;\R}�D�ׁ��N�iR\`�ϸ�%9]-��l`��و�,��ݹ�ր�J����C̭�u*&� UC�?� �B�Q�	^���*W`iZ���2r�|��/������p�Xk�GX�k]��u�w84���������H}���t)=��د����&��5�d$�����x�n�y��KA̡����$��^�!%s��=�Ǜ����@�U���%�D]���n��Pq-��?�)�I5�+n#;R���}�����!�=}�n��b�4br:'8y�̔�j�\L�w��G�M�)�$�T��U=;�L�9�"U�����iUI��Ϡ����W���:'��[�DEY�1p�&D��{CU��N]�I�G�cش�o���B}��o~v��6H&�%0�z��%�� (�����}�6~j�O���JH~�(	�o���X�=�F�`O.�8�����83;�����?�fnQitL\��I���3Mt�q�9p�L��mƁ6�:xj�G=f<ޕ�T���E��Ox���M�ݯ|K�lSa3w/��bd���m�ϧ����f>��.�H,�Y��e����j^�ڍu�ޥ6L�|w������:|�N�`{鸿C���"�⇦Fzؒ+)�m/�pvz�\�Ћ��UW�(�hgҎ�s���,�8z�1��@��F\jק['y��(��"i�?|����N�\��!B2�/���g�8��{�����G��n�� ���9^�"Հ��7!�p�.��*ξ$ ��T���W��9�3s�t"OB\����mj�.�(��Oz�շ�����9ϲ�0���0���S��SE�~���a�����x�}�)�П��=R����c�gđ\(��o�b^(NR��)�-���R
�mEױ���+��bZ~Z�!]�Ee*�쟮��["Y��{<���l �?m��Ƀ�UD>�4��;�@8S0�nYt��Lm�H
� n!�(�ɂ_�y�?ւXϊx���?�8G���M�˨�/i�lt)t>w#Q�z�?��T)�f������z��F��u��d����!t�6m�Ahr(g"�b���ڲ��n�C����0�R�s�J0V��bmX�o��B~+����r�V��z��4�p=Tk��W���~ޥ�6�c[��_����'�їw�"���7��̱=�-�C���zi�~�=$�;k�:�]{z(���Z������:�lb(�nT"��hE��eȯ��Ρ��;�:Ǹ�2X�x9�$G�`���=�y���&�r�P��](���2����Q�Ҭ��a8�7��}/�U�:�r��7��yܔ��_y���=���!���},�����CX�Gݢvd�W�?�~�ދ�w�	��X�-OL*�:�n�+��gG� S��#Yg���d��E8��4;��>�]��r�d���^��砀\>'m'�Io]��c�M<Uq��5�j���k�
R=%KHrd�3��l��$��@ʹ)i��D� �p��O.�-�j�K/��p|,׾VMj`���peR�Ly��J��Da����or_�wv�hB���d`��>�6��~����JvͨX�I�8P�
�0b��&�H@x�����y���V{��./����kz�\Bwb7`����F[׬�^�ێ�0 R���p+��?�&l@��u�W�Qך�w�>��f�����I�f�Y�L����O�#�wiڱG�?�T�F�2�$	��[�	e?肾�a��`�nh�B�,��7�"3��T�z�ё�Rc�P�)���JDI[h�U��7�,R�\��b;���:��@�}����̀���Sv���S��-����O�y�_��5Il���:u�u�q�',���,r���DQN�L�?a>�ދ>�f�웇�A�*�>,_n�@l�Q`��d����B�%$C��]���_9��T_��� � ���x��&|�Z�BZ�/�Ȏj=�eQ>W�{���y�"��s{|�u�_��7���n��Ѻ�#B�:DZ�}�� �ӌ6�L��&�S�����zm�=���&��{�4d��d���I	6� ��hF���>l�����(�	�+d���*��'Ǫ=���lb���5�	m5W�K7��Z�j�q�݌
�;��x��O{U���I�Ie�KL?�\��2��ल�DB@��3�Inx=0�y&��,����
�����^��;Q�ˬ̐B²���~���6M�B��R�kI)�
9�m)�|g�Q{��!C uwl���	ϛj��$��.�����3�ޕ����m�k?��Yr�B�h�|Uۆr  �f�<9�r�t	�4�RSD�T�u���jC∬�F��Ji1� ����_$�<c#���B/��͂�J�_:���m�w!�;�5��h-��P]"\��+׮�)���YȜ��9C;#Kn�Vr�E���]S7�1}Ւo�՟gp>�ᢾ����;
C�;}�&���E?�[��	�2Xt��14Y�I�_3��#ԥ�*�r*^��w�9��D��e@��Nn̏� ``�l�-��j_�5���jrfyk&Y�ݖ��Y@y��Υ���i)_�7���зp�B9�Ay�d07\���_�P�3�q������υ�Z�buݳ��Q�����.v����Y�~܁��a�k�� ^��E ʋ�D�mG�_k���o����˵e���L5�'R���jF���0zr)�íy���NX%/Ò���3�i���-"����nj̟�A��װ|&��TE ��oE�e���O6J�5��v573�FR��4��Qw&�^72�j`�z�kɰ����e���N9��<ʳ����S{
%r�g��ނja�w^��[p� pD8l�E�-�>��yZ4���	kb
��-��xI�k5mO��U�������w��%����P1��{�-X|?�\V�WwT~�u瘵p�ڨ�̍n[�O����������QmC@�e�s��9"?r��9��q��X� 3ή�D�{'�7��Z�j_�Z��*���KT����\z0�
>em���n���H
�5��o;p�E�TJ���
EP��)��/��S�#m	8�c���W��m%�h�Ggk��.��GF���A��#�ԁ�)�}�l���G�|؊&7�.�&��a�F�찀�z��J��X������*g�kұ!D�'�'ޖ2&2�I��q��1G�%�����JG6f���T�m$�Hj��������S����J֖�V(�S]^}e7(=�cn�76,��I��I��O��ӏM��dM�6��S]�]�}6R:�_ژ���$���b���ͥ~�[�o������pps0!x�`�����Q���_����E�3����
L�#��c��`��y�Bur5��ӫL��Q#Z�˵f�]��F� �|6���� ���Ɛ��֕��بt3���G]c│��v$Ƿ�դ���BO�T�o]���g���V��2��	5����J�;ߑ��'2Փ
Ф-<\�z�=�!�����7m^��'� ���I�*d�/�i&\�FL��m��"m�}y_�n�8g̳)<Ϋy�t�8F5A�1�
�=Y�^P�!@D"r`@��G��W��H�!^��h�P�X=`$�-��.��D�&�����5ᕴ^5��-ؗ:���F�U r�gE�C���A)hۤ��Z���5�5��L��B
OCHܢr��q�:��e������Ӫ�-��}{��<D���17Ԭ��~�Tj�f�lFv�����VF�,�����8�˫�`�VH�r�>q����p����<��G!P.w<�e3�,�X�8��F"�=�K�c�l5D:�����k��@�^�*.�1�q��!�KS�#��mZqyY�q3X+ɲ����W��w�nL�s�uC�HT|�˛*+��	r4�����G�boG�p|��m?e)my�-1�!pә���n�β³�Tn���A�"UlCm��>u�ϛn��:�Ժʫ�Jx �h{6Ԅ�y$��b��Rn8�y�����;`j�>��R\��q'�L�7wX�=�<@+n��S���
$9C��i5o�^�HS������n���S�P�M�R����2Pt��Jo�f�^�l�,GU�?�g����|��:�����~C[���c,�z����P��U��U5�'C �v�Rp��<�Ա㖳N�Y�_0�_j9@�� b�e*ה��%ի��B��󑋢l���C��;5E�E₌0��Xs������Խ�h��e^���NSAq�؆9U��lW�}���}��R�E�M_
,c��[��lSI��F�h��B�UW_��E'Q��rIV}�]o���->��A�8h��4��N���i�#���C��yF9�$�� ����g�R�؈߷ n:l���Nw�p����k"�/CV|�	���<ol1�:T���0&C��i�緣��y�X���� �v|l� ,�k=Ί�O'F���h㽦�����3�o����eΉ<��^ku��	1���jR��U�X�|���ia�q�6�:*�/���X������w_���OW�$!��Ɩ��T���1U�@�dLGaZ�{}#�ψ���s�~�����j�<i@��A��j��/3yn���.w��ά��]�7�n�/'Փc9_��,�oaXzC��l
>�%�k�m���+��3*�v�?�HG��m�OE��프�̖K�@Y��� �b6�B ��e$#,d3�EU�Ĩ��Ӣr��>��B�b	h3D��,�}`��g�K���$>�xEN�=�����������H�C��ؒ��J��dC!���66���>���ĜA\�Sh)�~�m�O� 	�K�)��_8��IT@Ň���Q��O�}	RxU̀�e�4��7V#~e�u�T \��%�U�W
�F�m�>Ed����3�x�^9�j��v�t�����h1��lu+V��*��U
���A5�F��j0���!R/%�Z��*|�ʋ�}=�K{z�\�-3̛���g�Ի8�(�h�K~]�I���GL�O�OÅ���U?�t�/�V���BA��:���g)��	�ZG��ɹ��2�P��S���U��ǫ��=[�ȘͰ	eEy=v���<�>��V����N�L�v�H@�Ƀ|�'LIPq�qX��Ylt��2����'̮��]Ј���
����+�w}LH�ƅz`xs��>�(�䲷�t�8�!w��V��9�7W�ҩ�/Plt�L���2��f(���+�0�-�"<[q��d���J�n�G�):[������2�<��b�����hE�Z���#�b�)j�K(U�@u�Vp�-�����I�f��+wm~���)B�V��+!Y�k���aܦ���Ά�����M٧�}�"����,�L��q��tC{�Q-�=Q�A�T��ވQ0��]��-l+u�7�|����+CiՌ���[؉�o|nK�?.pV�L�>T��OY$�NG�m���յ.�/� r�z��2��D%H�7}N.QZ��N�j'�o����	#c�+,�^������2b������w�9U�=����L� ]�4�7����N2��/-�M\ii�;Nu��.��{'ucƗ�O.����,!�-�a� �9(T��;��]Lx ����H��3���Bs�{t��6:���k�Tf�H6�O�d%�ډ�����qq��=���s�K!���G�e�y��VL��X����F�(�=��E�V�y!�`�9+��tLˎ��4H�b������� �"��ֆ�Pȼzd�C�ͻ�����<�0/��YN��d2�XÓhvNzZ�8Ϯ ��r�i;�%"	3,(k��L��I˖���^�7�O�?��i5#Q���LS���*�Ý&���C���	��>�?�^ d�m6',M�=��i����}*��)�U����8�
�s�Cń�d�=&��Zdk]TK�{�#�����H糆>��| ������{(-���n�b�RZ$|�53�G�i�ʠ%첰�[+��Z���N#T�x�7�5N��}2X�}lm��w��R7E���|�zh��/������1�\ۻ�׏�!T�V#����Q���f(.�b���� �����R���N ��'*�cK��!�H��w�m����RIX�	�m;�Uuk�u+>M��`-D�s�J��
�E�<��I`��b���@�m1��i+h.	6��z*� g�?�y߷%mE1>i�$=�ѱ�s4(���Ԛ�L���T�5T��Р�O�>H7`ˇ����y*+����L>�z�����	�!H����)�P?J��/lp<�Rb�:п�Fΰ��F6߾�T����� �,���w$�2�!�9��WL~u �d�ǰ�L�$8�qrMv���ҷ����J��a�ｂILy[�V�|
�fh���wCG�����'K?^@��	�y��:Z��Lí���b��7P�TY�V��"��2Ra����3j�}7���Ju���ԉ�q�-�3\�m�ڔ�ڒK�eE�fS����R\ZX�Q�Q�~ٻ��yV��}��Po�>8T4�l��Q�2�E22$��g��e���~�c�y��@d<
���hu��-� { %.����<��c8�V^�B=��8�<!`-��CO�C#����D��څ 5�X�}�S�L�i#A$�����PK�'ǣ�Y�gS�IUh���b���^�]x>)	7G*x�]����i�L�+d�Z�8��]@�p ��SoV8�'���WB�<M&�J�tQ���l�5V����W�X�����Db��C��)�W��J&���y���8h �T�4{w������RT�N��
�@��[XO�#���ˇ�L���F1��k�0#lB�v�;����Ϳŧ�!yxb����Dc9o���@]�@M��JM��Y_�����'^͆:��ЬS�=�#�ބ��%0�e��.��x���M�2(V�ž���##�
�QY	���8���+S6A�v���L~�Ro�@��Oi���sc{{j���`.�E����=1w��m8R���|�`� �ۆ�<)LA�*���@���(j��E��>��-�sP�|��+���6g�����~�'�G�0����G�c���I/K���cal*�qy�ҎTu�����P�\�J#\{��I�20�3�����1L��u)A)ݠ�JS?i��|4����<Z��1�u��;?��s����Ƈ2�Ƀ?g݅*���Z�Ʒ�35̃VV��ڈ��}.*bN��/��ah}�v/�'�4�" �0���M�%���{��݋F�*���CX���`���H�ҭF��U���p�le;�m�G���0���Z���k
��	�b'�R��I��|p�gs�4�8������8x�
��̋���Ѧ��(��=q�՞2��u��x��2����Y3��PY��� T�fQ�4��6���>�D��ݐ8���`7G#ٝ�|��
��_-��H��6�iͽ�<h���ZO��������i��36����s�9EtASudA/?�T��Ȑ��:��^��$:V^���B�8;�ˌ$�j�
�)��"j��g�㵘3��v�΢ZQ{h.���s����N {.HF&�*�	���,�s��{��Q�i��s]���+E���r�|'p�M��B��D.�^��ę�:�Y�4 �9U�VkbG���U)	�CRS��`i2{_rw5��!&5�؈h���!���N�T�^�wJ�tH��]�li9J͔b���R�D�j������J��E	�Rɿ���Aʹ�@�;�\�� ����J,����%%y�R���xEYjc��G\�X��f�S{0.I$	)5�0��v��F�
��Vl����D���؇�u�|V)��2^6
M�&w�tZ����Ш�P*j��mm ��Fx�W�C8��9=4��)Қ�t�g�7Wc��
�=�Ոi��N�U<�R-�_��Պ�4��6�,p�k�,@���3Ds���+�+��w��c˴�����R���ݮ-^Kn���ٕiq��cQ2e�;Qݝ��1#Yհ���2ԫ���b3b��C]�T��"at\I�?�Qb�B��t�鿡���2T��^�`�ت�,'���������g�Y+�N�$�=y�T�s9�	^s�,Z��?r?�<�$քT뮬��;��0��8��B�.?�0���e��mg�`[<{cՇ���b��B#��.���$�?QgA�Nٹ�g[�bE���Z��h��x���<���^�7��|RV�@2�Q�}t?�H�7^1d��L�ծ����,,��~��<}��lr�����Q��|G��LՀ��;j����ϯ`��^����ؕ�v��$�;���~��q΢�(���<F�a$�/�=Z^i �g,�9gst�eBr9?�G~
�g���o�Xܧ�A)�;>��:
�X����\#�X���`<���oqݥ��P5�IWq�����U<��2Z.��l!v��x��a��!��2��ND|����@á�ͣ�f��ƍ8l�0��"`��z��,�������h�9��F��õF��Dg��y�O_�������Ƭ�cG���w8_,fRn���I:���l\s! aQ�@�w�DY,�'3Xr���# �����/܋����r�.���
#Dȱ.Hk�y��5��-��#��^2�GMPڊ�W1Oe��-v���B#K�IP9��zP��N=y#�;�A��{3�,N��K���K����z�`�b���x.-�1���dէ9bPw���o�\�d��PB�@�oM0�l��
m�h��$lN�&��<YU������K�i���w�Prq�z��p��ⲾaL�RU`)Fs;�-Zx�Z�NN�2$9�)>8o�^�k.&���gyҮRjDjL䢲d�`�U���c ��X%u��^�(�`7��I:��?�v_<z��B]�hȱa,v���z*8�Q� �Ϥ�"�{q��g�TU��Xp���1���1�tsx�j���<k1�{������������W�舧:�o1�� 19M-��L>;u~�V�	����r�4�	Ҡ���~���5��^�#���^��F�g�;rØ��J�؆��8;��@yMw�W|(#�� ��E9r�Q�Z���	�.�ro��@5�h�D�e��O'�Ҋn��Lf���}��̵������<l���,qZa�l3��ƣ�-/,�ғ�+��u��(�odoQl .Nm�� ���؅b�s �ߔ�J�"�Hoe]�Q�k����j�Kk?�����l��w�h�8����B��c����4��0��(ΛXe��C�:�{��Tr��e�9�+Ց�P�2̩F,s��ښ�~��:�&��������p*�I[i�@��jV>�(�5�Go1d|KX�N�L�"��Ԗ�ʨμ,2(�xS|[�>��S\�f}^����pF� �z��p�׏n�@1�>��o���~������sIpa>ֻ��m�ӗ��R�̣ ����� �Hay`�]�2v-k?�t�(�vo��y}�_>f����Ͷ�ѵ�<�]T�[Y������ǱJ5��k}�s�
7[���M��h�?W'UJ5�	ؓ�l���Bۈe� j 6�\j�-�bo���wt��� �}U�yn�`l
���x@�c�jp�#�1-%�Pq0۬K�7I�%����y
��
���Q�hKc�O�k��Qce�8!U/�\�3G�&�v^g<%�,��ON"�#���V� -��=9� ��z�n���GG4%~*\c�A;֢����q�ǣ%(��]�4>�r2'��������G�+���ķ4TO<K�Z��굚�k�"֩���z�*0C@[5�*�O��TA���̫�]~��߂�?a%�"��+�yA���`�(���T��м��^~�`@����=����J��
�(�`:�ؽ,x�w���u�À��Z[E(N,�i��U!6"Aׄ�擥:>��o~0)�:�0���k�y�"�[} @�ڬ�o]��3s#PӇ��@{�2ٸ��p� Y�
y��"�r��k0���D�ܦa�_Uj�g�M�{g�b����g����O�%��,���'kZw �:W�Áe(�},VJ��}�����3rI#=��g���V�"�}�P���U���n�gK����X.�(�Cۺ����0g�I��IrԵq�\�e���|���Z��ꦱ�Sv�{z��"E���JFaC�Y���k
��qY-I���K��h�6��d��(U�K_7rp�e(�C�:!2F��og.�㉆�8�x"/��	�<.F���U�-;K�Bҭg�f_������cR;�ް!Eaì�tѢ矀.�F�!��֘Q+ �#$���U}	�#"�G	���Z�Rn.�f���K��)��7!9yG�y�ʺl��v.�r��7�!�q➚�P���i���/�3�l�^�&zN&�=]߁�������,6Y�F@@R�N�Z6 2�s�Ѫ������
.b6uQJ�d�$�f+:J$�*9 ��y"IБplt��y 9��0����A�s;ȷP��C~B?�ߑ`쏲�v��Q���D����b_�f
��ݻO��(�Qج9+Z��1��hS�=�5�[YBB����E����@�^�h3��
5N�jװ���k4�s��O0�l/��g��D�� �!��P� ����q���:��Ր�+O�v�t6=s~���'O�mG�i�s���� j@FZ�z�o�H��~Vʰ�]��]�^f��;�X���B�&�G��6�cZA������n2���y�oZ9�ˍ��(��F����`��1�_�y�$�q��[��` AF�����w,�W*�Zs~�
� G�B\��n��8�$AL�H�cI�/]"��4�xh���m�(�!�!x����<������j�B�[��t~��b�2�VYg+4����(�*	�1M#�D��Jb��݉rS$��7�7+e5Z��@~��V�/�`����jָ�J��zxL���]_Oߞ����{��"�?���<�}��z� ����)�#����W��2����t��T�>���(��'��<^W����������_+2b��� �"��������O��U}`o���x��� @�7L��� 'N�E�厙	��B���j�d��O�萜rq'��賡޶y[G��
�xB�yr\�>q#o��>:^�?�#�ɚ�,�oo*GQ_|�;�2pWo��b-��?�{W�DD:릡8�u7=8�x��f�⥆��/뫊�X'~CZ��A��������5�Vg�"/S'u�E����B���p`�e�uK�e�+r�[zseV|-\w0][O�]�i�D�8�����F$���g ��q�dIVK������G���opy��e�f��"z\v�ް�Q��C�q�,�[����خt/�<4��#;|b#��7N�T�����A1Z<8L�nYK_9|о;�Aua9#�%���;�m��8,;3\�w3\c_k�M��\e�&������Q9GM���K�:��7y��C�{k���T�+�3[�*,��Y�6�i�������ey,���~P�1^zM�B��N��D���iUC,��%�?�Gۖ�f��
�{��(������l�{�AY|�)&e�	�� J�#lk�؈�x����􇑭�?D*����A9���$/���j���#t.��҄_?~�t�(��d;����f́w[�ثP{��վ����U� "3�8Q��$z������v	���Y��ߒ�,����ȏj-ϓ�Tֿz�Se��T�
����H���� N�!?ʑ
�}�MfstS�f���츆��&���"�/ ��P�e��}_�X�U�-JQM��t@��!� 1��4��t HHto�t��$�K�;�nJ6��)��r]�3��A�n=� � ��d: �p��T�6�	o^[;�}j!���
�O��҆u�:I��-�jUw_��(	�@�\f��4BtU�����p���:r$`UNP��m�A��4�T���DPu1����ې"�AXbA�'�S/3�c�b�h�;�z�.V��	E�$�Q����*��H!6]*3w/B�{�W(���\t�^��c�u��ND!@�ٚ�ϓ:��AΏF����n�
���'2�ɋ�����s�d=���<�����e2�f s�ܱex@�K-o4?�t6�R]���$(�)�̜����*9��s�ј�>�U�X5V'G|Kb ;�r�JP���	w\:'&���ya�����U�>�s�.�9�n���KA���\.?�)B?��������{=��ؕ��X���z�wkH֬O59z�$�b��rY����l�#�4DY�����, }�j��f�3�
KsW#[0�B�ˋ���';��1�ha�3n���_� Q�S釞m�	��6d�ؘ_�c[o2!�^����9��b2R�-�J�s�~�n؁B�m/��9>�6ѐ��d�4k�����Љ�gXE�]�HX<�y{'8ϧ@0�mХ�*�y��j�G�T�8=g�qSR����(@
0TB1!E�������c�*��e��c�8i��Z�s��i�z �E�<�!Émdq�OW�?'�s�-�AO�U	NEr�F���/�}�J���Hζ�����n���yY+s���!���9�3=���Cd{̖P��78������n_`X_y���Jt��l����F��8�+Q�������%���ӄGb��~�ͧr�s��.	R�'�@�����Q�+���cH�<�b�N?��z
�Fh�\��!�I{x�m�񭞋����a�p$��*D
>#������#J��⮗l��룲�>W�zM�iZ�����U���yϝhx8exЉ-��=M4e��g�3���㹊sXխL���3�`�5n3�i���{_f@����a.���oF3>���k$�^7��J�H����x��.^,o��Q1U�<V�C��D��w��6�U�&�'�f���a��T� 3��gͼ��Q�,��2����u���u���f�y��l�ե$N(�H����n�-՜8��G�P�S&�ŷ쵧��fL��{�eN�-���g�Okx�q��x@]r8 |xy�3Ď�m�)6���l �M�\��7��&��`B�����}Lk�̼<�)��;*���c� xFH�U]��(�reP�l0����3� ����q�6�8k�I�t=Q,������p(z<�� ����RL0+��1��V��>�=݂R��2��D��K_V�P'P�T�Z�v9{��=����/�"DR���������,�A�ը>/
��̙�.�.���o�y�W��"b������G:~�&Yg�E� W��Wz.|/Ȫg��N���v��B_�@�9
�̻Dnw���;7�>H��`��r�g�Ne	6$ά���J+�
���1f���k�z��b�+Y�t�\F���K�R�`��%�U\�¯����d�u-�-����ʍ�Н�buE�9����a�xB��/��R�P�-c����Oc1�S�Ma�d ��Vۺ�^Ǐ���]K � q�s��Ք,
���Ԏ���r��`]���x�Ҕ���N��Y��.҉��⠠������PoE�B02G�\�.�ډ�)5y�Wa˕]��G
�\P����ȩ�V%���N�_�FB&)t�r�*QF���Ӧy�<�;���a�~��_�:��S<����4��/�n������Y��d��K_��a��VȊ�Q(w���ݲ�D!�5jS��M��&��Z�b��*���m������s�LGr�heU�o,x��[<��I�p�w5a�-K�p	�C�u���tfd�"Q���5���V_i�34��U���Ɍ�h�����/�ɭ�(��q�g�a����1��sb-ܞ6�L�0�ZdgR�l�!��Ld�,L$�lo̢�1�6z�3GkbL^G�@��e�����>��!��X��o]Q��d:ޕu��i*2��M�3'��8�PBlV#LZ��D���{�)��D�����U��(�h|����n$�����`E�eڞ�I����4W^v@t��q��	���)*���N̡Ĳ����P@��]�X������ϳGU�F�8qd3?�K'ΙA��^�<!�+������� ��Je=�󐁕�
����z
ľ:�rd���/���x���O#\��SN,B�݋r���Ӷ�����I'��	�W� <[�P+�����_|ܘ��B�W�Y�D�T���S���_��M�U�
�=�0��<Y�:��w�A����ȩA�W�[�Q^]�[?�[���1�ע���'2�ꃱ�߸R�C�Й��(�KG汲���:��i��ÿq��gy�i�.���2)8�����i�
;s��_��}�	lp��}<)��vD����6�ծ��/�٠��#E�IG�P�� {D[V�+�/�Qh�P�ϭr ��e�"�S��(�~��-G�zO���dp���U>p�9��mr����������d�vTP�8�O|�އ�	in���qZ�אָ��I���*��N�� 5ap?�ߗ�����j �0�#�������7r�P����Ȏ�_�	B>b��>aܨ�w�������i>�����n�{0�$L)nL���ӄ4ھv�Sz�=.�(�2a�����CuΚu���Hd�M��6:%�����wf*����.�%���y��1=
�'**!F[�H�@N���DL�{Z��|��{��t��_=쟷�	Z��JjޥO!���5�pv�*!�5�L�[q��M�8���Z/���N�riY�jZ�T0�{�B_J�F���U(�y��M���Mj�����^�/w�%��$|�ل*Iɷ�z��1�kzc�C�]l�����OyO���z��&��a��_�z��Ԑ�c]�&�z���=�o��ѳ�˝8K�}�5i��DOi�I��� � @��׾���2���"�9���9���׈ޓ�ޫ�L~��,o��<F)�hWO���%WC F���{�.'���@����
��L���ꑪyj�:��} �O��rm�x���]:W�ˑ��u����.ٟ�\T����1Y\0���\�*h�U��l�S��$W=yd�k�]ħ��c�����5��!�k�[c������S�27�#ҕ�e 7�U�����Mm�0;�r�����J�o}]�G�ޱ�$�@�|gYF��U5��g,0�{��Ex�3�6s��M�K��0Ka��ZՆ}x4�]t;'�@q��XI@�m[��h�a�k�s�+G�L�=�����e�zo_����rh"��6�GdxP�r����}�~c�vru���.���ߜ�e�31��sB���~~����6��������^O����I_X�-�D^.�z�d{,���E����I�x+���yj�j2�l<j��z
��:���C�u�l��G�!Չ���0���V�<ɬ�_j�y�]vL��.H]����lf���J�V��x��;�'!T��Ą�fIA�d��쓕���1u�z?l�[<��:��;@l_�{{�jYw��-&Syq�`O�B̝	M�Ԗ��צ��Œ�W��HqD��U���!�*e���U�v�cԲZ}���e�JrꜼ��^LY"y_�$����c۱��ax��n��jH��F��V�k<��a����iᒼ�����ƻ�vz�4_,�e~�8R�-���]ُR����qu�M.$�>��y�~\�B���h��R �o`Q,��X�?� ��1�҉�k��5ymxa�wd2���N���[�ߘ zT��Y��'AƄ}���|,Sp��v���[?�O
�J��d��-�t�����;x�"����Y �Csjx�$�x��Yb��,�D.|V�5Rt�z�&�|��&��A2�o{9쏚2,� ����Y�(�M(8�p����H��=���q1!����,�y��@�,G�V<��s�j�7����t1���J5-��$��^������B�}_�\��(���yzB$�Z�;�����Ց\A#��Q��R{{��u�->��C��5Y8���0�~|s�ͪ�{����.=�._�2�w��E̑�!Z����-�=�/��(�B��f	*��Z��8�!��ݿ�{l��+��H�����3���0�v���v�r�U��*�,�9./�^�zZ���z��������Ǡ���ٱ.���!���cxω�;��or\g��
�{�:��I� z��.��d3��Sؓ��Rs��< ��%�7.'�QO]{�T����殭*���y��82[\^����t	�3x�t�wU�^K�j0��Ċ<��41�1����s�T�V����?p���].��~	��cS(RMl՛��J����x��{�z¼В��y��?iI�}�J2����R 7Ռ���y@�I��߯c�˦?Oe���(p)xx��|��Z���TX�lז0�$F8P`�dg�CzC>��
l����1��ɵ���P,�b�IJ�q��,Y���B�hLYt�_��[BZ�M���"��Ը4,����a��R�6�m�t`���}E���X�wChz�Io��S�l,�z:�m�Q��-#��U��;�G�p�*x�~�>��8V�H�?����)516������}u�g�~OÕ'p��w�~��D�s���9j�H����Z�+�%�H�;/J�%��r�|�e�c9/�SY_q�Me���;��G֌&��`{���r^�e�!�u�
�}&O��20
�����d�IF�<#e'��F�u���3�Df+V��m��%���h�x;��\w8��!��ȍ7b�J�u ���.�\P*�ΝC��[[l][e��k�-�%��/]v@�V�߶8��(�n��P�[��_����.���4�B�zǕ�U�0�qr�_�32�q�Ua�}�1T��P{d]L>���%�����ά�C#L��̓n,��Ʋ�UT���k�J������:�਱{{+M��|��l=�-~�j�9�|Tɥh��+��F<�i��{��(?`V܀�����sd���*.�<|��"� �����e�+���I���Jw�5�<�@�R�
4��
�L3-�T;��sET��]y�(��w��+-(c^�_i܈{g�:*��S�{�(;:cH>8�?{,��e�����o����s;<�6B#�¿V3�CZ��������P��oJ`,�կ��_�NĶw�v`�&���r�
J�O=�`�m���B��c�ۛ)�p���W�]q��s����:��8�?�lX檧J�#b���g�����C�Ƒk]l�x*�J,�칢�����ލ�#>1ߋ�V�Z	X77����\=@/=
�ZV�?�$P�7l���e����"�|B��oܭ(,?so�!���a��M���9P�Hz��"�L)�1(��v��_�)F;���YN����C�����_Z?���zy%p�[�x�-y�%���uXų�H4��ȑu��ԭ��T�㛗�s �22"3����%�g))�OY�0ޥ�6��^`��F%b��/a	�\��$��O}=�XN�UJ.��ާ�+�NU���P��=,·�Ow�����g)�u�^Q�
K�<E�j��?F������'��~Z��~.
�ڲ�[� �m0=m�.�U�H�|��X����Oik���d۽�%'JY���Q��B�c;�m�`���u��Pش�@��2S��gqj��PÞ4�r�5?���}��{���A�	5� �~ѿ�B}��!�ߕ���z�W�Q'�X�C%��폨�\"��{��v���N��{f�OܲV�h��FU#<��nZ�!�#OI}�Cֱd� L 6�܌���܂}X�7o�g�ubi��%��k}�˅��O�L�p�.l9���l`��=e�I����}���f�Ik�����F�Hօ,��}��_fѓ^��0$f=G\6��#־��!<���Yd����(C)@�W��T����>�?Gʫ�W���)�F��V��7��$��$�	7�)�'Z%[uhH2�e��Ҟ
��W��ۖ�����Ѿ@�k���R��T��t5�,���$��.r��>SN�� _���C�G����A��{7H��'&�B��P4eW�<߷���0�}Yb�V��R "�(��pt��=k:���!�3 ��L�U��*�.��������jf^�¬� B�q7��B<����ˢ���f&�BC9�I�$۴�$up�Y��ƿJ%�<DR���/*�Ӏ�w�%"�3Z�|W��_Y�츗X�1C��Jy���|}9z;�,�+�4/g��D�n�~�s&ـ�q�=m�"w�[Fcb��η��<�������y�4�Lϥ�����Ӄ�}֒�]�>3��!�H��T����-zvlK��>�9&���e� V�e��V|��*�"2����y�=�WIC2�|\����f�d^A���hxn��z���E��X�(1�c�o@���#z����~�C�pn.��v���}�V�C!9�\v%�Eb�ͦ�ID�oԸ�$��2�/~��ZHn�*�+��|�*@��б�����˫���
B�n��9�c	���R�!�IH�>��\�Ώ�d����������5�E8[Sj4z��N8���i2��]�'��<�����4��8�q:|<h�����/�?Ym�G"ۖ��z��A�j��ؑ�}�����kR��n�rP]�i�rK�6RN����t�Zp0,T��se�!2U_�VO��k#K��P�ۗ�A*:��q�]�u���HE�����r�Ƭ������E���,v���Z�/�0�r�gI�J:H皋u"��L���=�#c�i^���������g���.ȝJ�A��#Y�aU�$�Eg�:���y�{�߷���m�=�0�!v��i�ɮ+5̜Qc�Ţc6��)��2��"�B����Q(���zTƑ}� �Yg!�ay�%E��2�n��0�bDi� P
o���7��u���L�K�������sQ�#��w��a�f'����	�՘�,&��H`P��l���ðd+,%�B�����l����o�<�(���/�P�Et��b$8���*�pEq� ���"�?V&����]�M����
��m�������݉�^��A;�ŵ�e�*���� Y�j���۪��]�s/�߈�F�I�r��z��\�����S��F+�!�	�3�}���� �Y��*E*�&--Y�D:��&�Cԟ��E+y9�p��!C1N�����HmG�:v~�=���Q`q9�[ -(4xu�������O+����;)��ں|�ٶ����4`֕ɂ"�O"�Uw
�30l�J���baD6D^uM�]��?���I��A�������'y��W����� 0�%�O�`�jv�+s>�Th�ݖռ�t��)� �ub�q�ܢ``����jZ�/v��b���O���74M�o��e�WI^�
H�D���ܘ�@r��zä``|�eG~���M�H�Q^��m&���͸�z�&��N��;��҇q�AJ$���F�u��]Ð5N9*�5�yΏXe��5���#t���ls:���2.��.�ţPU�Tg�]b+=|y84��/_�p�k_)�R��T�p0p�iC�o������b�G�҅��F�&I�о*x�����~[������M*p�Ifw{��X1S��r�0�.n4"���X-��D����fU�F�jzl�x{��s�� ������Dhﳇ\�|7�7r|C��W�j��
�cQ���rnw#�`�b_`�<���֮����=(�'�����S���S��0*����G�&O}����A+^B��SΟ�b����v����z�jC��\mr}n�{6�~:�0'$g�v����d��[������G�岮�Xy�nP��o�w�#\�1�	��u<�u���)|˫@���`�ޏN���S�o4��Ö{����CCXg�p$���p��T�� ��X��bv�O��y��u(��ج�\������vI��o�i�((�{��Bc?U�yx.l]�=Ͳ���u�M���j�RA� =j�r���TtX�Ǉ�7�į3�����c��Ј|��D�=��w vɭɩ��3��%�s3�|[�g�xj�1�>�����iC@N�<q�5h^۰��zԘ���h��6JQ������K���&�/�b���=?~*f�׈eXv��
�T�
j[��4����j_Ey�u�ڌ��~��lj߹��rd%�R��y�B�=��G_�J?�2w��x�ul����K��Pm��p6�A�G�fzO��$Wu�1�T���?��������*�c���t^��c�C;���rDEU���I�Kl�ue@��\��u��A&��1�{�!0��5��v�m��& >�x$N

M��W2u�$U�3�+s]�_���r��[�u@8p|���j�~�Y:��Ko;�s-&�BY�|@�8\�%�@���E��q�M�R�D?�Ü��ٝ:��M��7^�M���� ɛ1ә�T[�� %,����\�7��n�f��#����X��T�������d��w<2��I�TBfK�HY!�տ�5w(��υߣ/Z!(���L;SK�Z����h�Ƕ��!e.��m������
��'`�x҇��^�W�,�� �_KUف��2�H�6�����xn��/��JP)��9ຈ�p0���t����=�I�YL��$�da�^�!A`س��?���}��js�h�b�����;�=����|$DF���s��脭D�	�S�[�aZS�2+�"R@��<��F�P[�!d4���L7�C*f�&vO�7�����Mc��=J)=���pK#X�L�-�v�Ȏ�k�Jm?`�N Q�}F5��N?��[ȗ��5B�A����evc9�ߢo�;���'�X���}NP�� �T}ءb�2�ë���=������)�Ι'���������<���t8�L�5"��J��G��!�N��:��<������kt�X�c�O��W&߃���ۉ�h{*�qxP�:�`�:$���}&iͣ1��58Xu�s��P�;��w��fftB�b�ti�.na*K�5��	����>j0�����5u�yv�N�4��.�G`��^Sw�aD�Y��u�9�L�~�35Xq�c�M�p��6ЃV��'T�!M�Ngp����������Igh�� ����/Tr#mH�+ �8Ro���e�d{�~�SU���Ёi��ee��b�f�t����{�M��� 	�=�����F��M��;�QP����]��P���p9���.�[!������_�2r,��jbXt'��u�B�r1N^�[5��m\ƥ��L�L��?�F�:XS�;�O	r2k���ݔ|��(~��ʛ}xOvlݲ�|D���	!���^��F��D*KoZ���2���&&%l�逰�oI��-P��0�'��a�
�P�"�7%��G��5�!� ��$ї�S�#��@�3���YY޽��fO��֩�:)}�9W�u螰D̞��Kx�Η&��I�s~�3.��!l �X�X��;ŸA�3=�t��|qT�y��ۄ ��Ň����!N�yn�!�N���UH��{EU����c�L���9Xs+�k;��;��_��
II$���P�U�Q�H%�J²o<d�]r�K$L�Sk`�7d�������Lp7#x��=�E�d�Bv�c��|4�D�aJ;��@�`%�Z�lJ���`�[$�d��w�~ײ���m
D}�!���1�w%좍+9T�v�
*�&�3�X���G�[�u
.`,9��f��;��
��������A�&����O_�T���c^�����j�M�n��E_�-��F��-'���i�M���i���>2t��P�T�GN�g�؄�o�P+�#�y\��5���w۸.��Ik1Ɉ`$[�*4y�Rp��n��YX07U�{;�D�&{�*<6��^\ĝ�IZW���?v��v�RZ�h�P���������>��|�O�Y���2�!��ޑ�o&��Ӑ M�N����Y���)'�p�}(v���g�?����З]E=_���H3Ig%�,�!:��f��M���Oy>z����w�*�F�4�aYG'� �]L��i��ZWB�@�&�'QF������p�uj�@[5�'D\Wa�'�Xh ��v����~����_P�bɁ\p�Q�)�P��s6��c��N����~����r<8j�Mn�cʒ�i%`���#�aC����=s*,r��#��j���	�Y��Mp�@99�d�����k3�1�(.~ zf`i�~���HG�+���P0!���ꋬ��u�]��r�j\��t��\�����<T5z��H$|9���t`Qٝ���I$-{���z�|��ߠ��
i3{�hCٺ3o|j�*>��lOM6Т�K����c裡�]z����@UtUHH�?���`P�J̊�Ѥ
�w�j�����A��ndn}��5�M�Hn¯�M��!����S���/�����W����������X���y����ۜ����4�� ���6����+MG�<=�:�W}�Ô�bj��_���҈1@������o�rM�]��	?�w�8�oI4���]��h��o{�!����&�F�ĭ�$�xPS�Nz47�	k\s�-��q
�m��!qp���̙��|��7+2�A��=� Fi;W����9��y~������g��	#�n8S@�=oo;Px���9�̢��O�Q��KeJe *lI�a�#����l�3�/�o��HQr��|�]��wL|�����4^�E�N�D+�i��Y����r�q�%Z�7!�_����ï���nO���ׇ��J�2(�����n��_���a2K���X�����Fm�?ar�{��,���ü	���Iq���B��K:7�Ǘ�s=ՙs�&A%�ۀ)��9V�b��7��y^pr�d����"�e�����y A���J�H��&���3dn�U��O�����I�2�~��>k��.��U�������ߊfıh����\�K�� �E=eS
WbVCՊSBB-��_�����"7�V�b�-�L�������l]�8�&DdH�e
e/��N;��ԃ���DJ�b�d@� �l����_��	�xv����� ��߃�1��&@�B�tXM���V|-�>d$�`�a��^u,�+��q�uƴй�������,6|$57����G!]�%H��bv_���`��/�ۏ𦰥�g�Z�>�۬��u��9�� �r�����\�!�������bU�)\�M�y�ߌSc�Vnp̙?����`g���i������'�0�(��6�b��#���߿f��6b���̒���,Y�u�2,��q �t�uA ��P�J��":.�IgnI����T^cZC�7ȃ2(�W�/�]�Fa?����#t�
���g���t6�9T���1ug�%i��w^�?��l�sY��/�4p� �Xn�1a!���y�+�FRҩ��%f��70Y��W��ԣрYle,�loF�qB�i���gTw�W�-��U6Zg[��4�zz��_&F(e��-�t�׌O�ד���v�����'������W7q�0ˢ�[����e�	�¾�;\W�T ��F�f�a#�|?I�L�]�3)]3dđzɈ��o{���"��~�f/|�4��C���{y��Yt��2H�@���b�| �CQ]1��F��vN�	������h\h�*�]�O����>�ncaֈ�� Jv���&}&�<�GehP�����鿅n���Dc�|l�E!��.����!�(R�8�(�����m3U��7:/5�䮘-�ABAZg���ecj,z��F��=�q��)�D��a�Ǧ�|�J%R�*N/��K�j^�c�����s5��>mN�];&�W��+�B�Ǵ��g����7pĪ؜A	o:��fI擐:�p+R4�Im�w��%�Q��VBI�t��?��+������S͘�קT���:�(����ݿ�T=/��fx���YUI�[�a匆��줘|n��@��I�Ը�C���Ӯ�̷t��Vs<A��y�tz&M5��� �i���t�=#��{u꾓;E�4,�;�ir��*�?�ݐ��	C:�G�[wp()s�y�b�P,ڪ�1���#X=�� 0eŘ/K:��e��]�-fM�JҼhE!o?�Z���<�h��"��!���7W|�m{�-`�+$i�=i�RU78��Pų,k��0h�_��#3��&�B�t�d�)�>UQ���[�Vzzh��왖�=�+�ڹ��?R���A�/s���߻��� ����{���a����<g��BCt���r��_h�[��P���fVᕻ���؊�5�>��h�I�p�>�Ÿ�R%^���b<<��AJ�:���5�����������䊾���_�2����>e���՜j	��D-�9Pl�	<d殻�����#��s��d.A�WX� <Y9�|6��N�9� �W��k���f�����N��;���E%�8��"\ԩ8�v�c��֯��m��A�x����.�Za�l�"�R@T�q ���$�.5R
<�H�!��t��o�r�c�ʹ���{.&���;��,��a$/�P4��_�֞>�d�̏�*�^���Z�I/#-Ds��8f,D��rn�b��Ҫ���6��7O�p�A��ڙi�*�P�.%k���%q�e¶�gp�<�#u�aW���ϣCDI0�SC�DT$�:����	:�4��͐��O�u�C��+��.G��V

�=�(wF�H� � ǋ�<�PPp�l�?��ZǞ�v_��=r�<��|>���Ds����=��X��`#)�dώ?@%�J (�)�%��g)�g��C{W��ǰ@ڲqQ�b�
��6�Ac��LI5*���6�&!�E�_�qv���p��Ѹ���P�)~������}^i�3�h&�T���$�G�bb��f�tSy�%��,!���t}aC�&��"/�4�;����Uv�y	�V�K�r�A�ہ�ԫ��2˳�$1�g ����<Cl.0�.0��f���z��{��J�TR�C�x{/r}p��D�,?^\�F_G0��<��i��JI�T�`����E>��׳�Ѓ Q�oyr����u������ysne��SW�O�'�jR$#�U����;��{��]�Fv����}P�T`�9G����B��Is�Sb��4�=���+�=���'5GU�{�������aҩ�	:��Y��:�M�!���=�%�IFJ (BLj�C�;��)m���Γ6�d�+U�
/�]�����A��O�P��S���9��*�|']ω2��ѝ���s����d?"'o�|8-W�8���[��i�����N�tSޯ>P&9ת��O4)�z-���d\1uK�S�\]<�����z��KEųSd�R��\+�{r=�
�R�@�n������s}��?s[M�{��&A�͌a4)���
ꤼ'FI�x9i����0	E4�X��EG4�@q�~b%��>��`��<{�K�����1bì2�}�xԜ�b��
��ie� E�䛋�
�x��_Fk4��j��)���,�;)M	v���������t���Xny����l�rR��)�/��$�P�9s -�+m��\�ɽ���lB���Dt�*X�]��0f��r�'ƿs�7��*� �!��"F~OΕ��Ƃ?�EB1��i�� ���=h�>�E
Ɗ&���cZ\q�u弝���i�$CB�d��ķ��$�^���-T*�$y
���Pi+���0o�GK� �Ŝ�6L�3��O۟0��t$���E��LL,�T��G�i,�[����?1��5���Z%\]�-$���T�jϦ1�[�����~�r	��E��K�O[���3.�Q`д���6g��~c!���W����ѩ�C�K��JFY�v����&3;4[���3��v�� �a��/+d�i�Wꩈ�|d,E�u�Gn��U�	�g��(L*�<�!'ղ֨в&�#��o}	�e��:�9��w��Ne�~�$�bYt����Zu{u��я2�ض��cMq�2W�����l�̒3?�?�a�~K+i��׽8)[�֛ʃ��Eѣ���;/FE�L��z�?l�*����Ⱥ�O_�\4���F��P�?Iv��B�mƿ=r�ޕ����FBiv�őM�쟄�=��e?�mG���[���ƅRT��a�P?]�y�㸵���u9o�d��6���㌃�e�:uIQB����B��yܵ{�d
i��Ga%0$�I��xK�%6d:��5��m>i&��̈R��]��CV�B/��|ܣw��9��g���^��R[F�E���)Jڲ`��+��'�/��ٖ�b������gAe�Т��dvV�l,�x�%��@���.lI�X�}C�E���W0J�d�V�������&�I_E��	�@��1��ŷ��Iu6�z� ��Ǵn@�xi~��:%����t9��%n�9-�uK�D��ao|�1ձ� 0��V��-�m�����=Z��
���{n�Br}���`��_�GZt��	t+d(n{�}6�
=FT� �����u6���08���'�d���?�tp����z./{3�(�S�L��^+�9��y\�׌�j�3J�m��?�Oвi��HUD����P�9Y���y�!W���ה�2�H�H�����:5��+�'��uh�z���o-�"j�ݕJ�bb�FgZ�-�v�::xU��n_4tc�Ԡ��&g��Y:=��'�"��D:�)j��/�Κ��]t��d=�'\���,��k3%ȳ�C��R��e��04/���2}���1V�zA�mh��2��^6$ǩ~'�hn<������̊vČ�F;��"Ȁ$����Xg�Q�%"[��A
G��a�3�,D�_�ѯY��1��R6�ؼ�;��8��]Ŋws�x	]�*��Z�rr������X��U�S����k?�iCSp*�ʼ�N��m�ˇ����Ʒ:����r��/���N�����J��q<�\@D�{�;�G	������f����0�5J�-j��p���&��̴<S
��4�3'i^R3E���2�2A���9�F�I[�k�Ls�;Ek"���A�_����Y�"�WԛP���ZQ�>r���k:}͔�lCn� �z�H?աp��a]��(�)1݇�Z�[����9L(�٪f�^�k�v������3��k�}ѠI������QQ�
e|{�J]l0�s��-Ǡۙð�|̹כr�p�����I΁��\�������<`���$��G�zfZ��(�Z4qN��I�u`V�,g��R��é�/'��|�Ň�Bf�@���"�.о��\KoޡE46xУv�ux�+�J�w�T@�/�߹M�S�0Y���/��S|�gυʝy�Z$�"2L�2*\��������o-������L���> 

�a������u�o��r�n<p&Pr�{du/�� �7E�=d��&^���� $7�!�m��n�Y��:s�Z7	E��+i�Ό�_�,���Y:�6��Hu}ũW>���%1dh�ڕG��7���\:\d9a��5	�i@v,k��h	9a �s��Tz�3���ޞ��?��Z^o�����^���  ~+�d�5.7��7>!��ȏ�h�j��^�~�$ ?�mL��d��`T��B�T�Yp�O�+�)Fy������`"P��%6i�Ia�@�x=��D�?8��=�&<���	��RYS2N�l٣!��{�,ڦ���e��f����2S��S�po�Ġ砕�k�g,��Q�ig]8
,2ɟ�cyN��i(��-^$Ö"J�&��l��Hos��g5�%��I�	���O���	ڦ��u�YaFZ��T�Wa9���H���gv�� C׸j4��ʯ������~�"�<�0S�#"O�X���fWn�������;{sXRZ��H���G��E덋o�E���s��_:�r
�W;�8/"S̬^V��]&����U$��(21>��fa�W�`~�G�T<ّY��%fRr �:4yN�\�ϊ"�����%�BD ��F�%�������y�^RV����^�B]v|�
0�h�ÿ���/��=��JW�ƀ���I�L(�Oeh�	��o���	�8���K@�&�e���z���"���z���>m^\db/���B��pCd�NoX�_|���b.Ҙ�̼�vQ=�H�4�|��Tޝ#a���I�U7�DJ�#�Q�W;;j;on��ȉ�F�|f&Oqxq-�^-�/���F������:��L�f�X�8/�#z	@Y⭩���\�eDS�31���Z5[�pA�[)�*���4u2�2"�
��і�~�Q�@25�Vp�ʣfU��~g��6�ل�Sz���o��3�o\n	Z0�g��=lb��u�)#a�%��!�\���Ds�'2��^xѩJ�[�
�Py3؆���<�t6����-4�M�}(�E*�5$��7M�HL����͈f��Y3$4�n^���7k�����V�t�L���<�ϲ�'��J3.�/��]G��8N;����A��$y�� _%1��u�j�^�b�);:���2�[U�|���a}��@�)�.����Xe�����bb�kq�)�]�G6���ռ�7ya�.=V���� D�	�����X2t���f��� �a����\mdN�9�����A��C1������z�n̴���$w?�����~���Ѻ�h��l>2]$�Q���=��o����nJ�o�o}��B%օmG�ej���7)o
�GM��*�����!�c+�o��z>�̳&� ��L���:���J���4�"9u�1��9Fͧ�pN��d�a$��hHIbp2vz���"��1#���]�����%S(�i�馿�����/a�b�l>�Χ�&�y��#Aa�A��+���n�V�;	���X�i^��j@_z4��^u�_Ȃ���+�^5���9Lĺ��o$AQ0~��=�?�p�͛T����`�<�=~�����WV�Pb/S�A}�L{�P��!|�;�ȶ�>�A1��M��m�e^Z;�D�)��ċ!$�A���*�1;�3���Z������8��4:��|�.daIR]����k�pю��;�K����y8^��LS-l�Y(ί�0���Çr��tI���V��⎼���ꃋ���˪ï�4T5t'�b|#/�IH�@Q���;?6�k�p�����|�8>p�l��+���#Ʒ�KW���k�^MK'��������d�f��bP�1B��,�v�N`[IauGb{���	����ˊT�)���I5[�&�l��'��3z}T
<��q�LlwF�[�A�#�Cٺ����1_dj�J�����f�p��S�Ч��ԢC� �x�}5�[S���~L��(�����i��c<�؈̛�	����{U�����/�u�g.�������O����d�C�Yd�^XS�1��]+7�E�Lߛy0B�P��N[(��q�� `6��.,G���*1ޱ{��f��e\q�S�����uд�D���e\GF���a4� ����Y��l5��w�	��L4}V^���V|�A8�1T��b�V����S�>�.`�١�%.�^>�(�Bc"�\��	n�p�	�W|���X�d>�J&I����`ן��ư-�Ҕ	�z��J\��7���޷ն���6֚>�W�oH� �4gde)�B��BqK�u?i���F�
a�v`��p6��ς:OȐ�K�?��?Z1%̃����o9��9:`~LBF-�4)e�!�����z��џM<M:��V�=�#.f�(�Nx�	���~t��l;=ywt�2�=��R֊�!mm)�
��qF��ɞ���d����@�0���6>3gR�����s����ȷ
�r�Y�yI�������-.+R�8l--V��.�"�]A���WНe�[�)��F7m���n75��c,�'`�����I5�>R����H:�w;Ɗz�J�-�����8:t��E���Ӆ4��A�)H�Jz�+����p�� 4��е�,�����^$�yM�)WB��<��4UGn�����L�g��i꼜��n�b�ʾ�i'G�ՍN�~=�m���7�����-,/KqF���rQ�W^&a�L$��8���,�b�-�v���ȍk����}p�ߧ�Cj3,����]�REE� �kq��TƵo!pS�XmW4�6�x��rO�a�g��A)�i�wL���P�!uI����P��ܕf�3���G5�G@��k�֗S�GX��SyՅl�pɥ���I��Fj�<�i�%�7 �s�I�z�؎�1��f?/I��
,J���Mܵ���7E�uT�]�<�پ��o)@��pz�w�ۆ~%��@��nN�}~����v��T�e�I���}�6�$]�r�ߏ�W�Y��3�k���p�>�i��໶�b-��o�-���Y� `��y3?����� fqϬ�a���s��ɣLw,\1�/XSl����r�8��Q�%�ME̸���?�HW�Gx��{	��6�N ��~� (#�0���An��?�j�O�%vO�=^�B�B@_g��
��m� �x�[�|��Q{�Ð)Yvآ5p�Z8%��v�Ր;�D���kv쳵����� ���^M��-����.e�CՌ�È�/GC�(�62�u�D�}�_qX���fο\,$r0�ԀcҡJB�bd�[�x{]?����������j�o���+U<�`ȒMh�8���	�.�J�p��KL�4�3&~9FZZ�D�s��8j�H�k*�o��\��6Il������,ui�\l�ߛ�wlxǇ����W������1!���g�4�imzB$��vZ̤@�*T"�$U���$<�`�<����.���m����ir��2��$`	��E����	���r<�g���<s#yI��t)iy=����R��b��#�/��Tcg��$3	2��0�B�v���S?��A��#�!a<F⪄L��T��i�Ƒ����HtЪ��2�=<��r�?����)W���:�6��)0���(�S�]��[�{=��x��l	=�d�}��M�`eW�w�\d�9�=MR|~\�W��7 ��;��t
����
����N��a�y3Ng�˶a	�����l��C���if��!c��f���=P�ʵ*�q�J9u����;��n/�G�|p��Q���cF��t����on�:q���:�����G�~m,=����������w2{XL՚�鴅� U��f ����}���6��Z0��4t)F�\�h�3�Q=�>Mp-0ma��^j�%W��D
5�gr�g����i� �p�;�&����\��-�q����k�\l�. qt��NÇ�h�"Hd�r��O�V�+(/ d�5��ڃ�K�j9�
Z�g��bU��=�h��.8�yhj�{\:��N�@�x�J�����׿�@�������,�0�gh��M��W��$w��y���+˿�/�c]�E�X�=q�a�4*�K�ۯw�hu*, b,RH̓�)%��>Q��LP[u
?����e]R8E��>GPr�ġL���|��Q���ŋx�������B���*�K{�.����5sR���.���7��:��?�ae��e�!Ak��m'f�u�i���wp^�%7�R'{O����/I������>V�z~>�kL�O{��X����v�!m�Jn��'$��S�Nb����I�dnA�f1��؟f-}<d\�♨Ae�A���8�q$�qT��d�a�U�f�#Ej���%�>;��۝X�Y��S]����|�#3�����stu u�S�d:�(˸~�G�UBs�c���ő�	7�F�ykc�
�Ð0�ǭ�E��yY��W����ˑ-,�&�	�V0p��K�]9�%-�Y�u"�b�yf��j5�4�[�9���@=�z z��'��iC���e��D����Y�Hܿ	[�d}y��F� �]�r�Gqx�"�YO@���p�˸��t� A� �&*$=HzH��6V�0N:\U��[/���ɮ��7����r:[����Fl̗�L.��d����dޏ��9ތ_�s���D�[/0S�1 1��(TOb��2������݃D��Ƃ�1Kv���x���	��9:���o�s���Y�f��K�����2n�3��{�A�H����ct`�Hdm-3������?����L�w�������ʞ�L-L�mm��/���sH. ��@���q	i/W=}H�k<jP~NEKw�L�"���Y�3��ƆC��^9� �Z8r)N�Dx��uv�y�>B�m�a�7�e��A���jv�T���."J��k�au�j�u˰!�X�/�׋�j�������7�,�o��*�o�80s��Wqq<�L�P���S��g?���ƈkWo��R�8�jeGh�٢���h�@�hc����S�.zO+*y�������5��9����a%�Rb�Q��_���f.Sy�W��XsL�H�l�dPIBu��z��oH[���n�̌��ji�°읐"�͓�a�S��O�T��X���)�H�&'���6^&�{T��f��X������j�����[n�:+1\�5���?~�CA{I$$���bL�/O�������.4��|P��.i�V^Vf5�H\�hs^��$Q�u�'xH	�՘6t�j�,�����}@�S_��׍_���Kx�]8�1�1��D�}JU��^�ǜ�ͷ��qS�V�7��iUt���B��6{Yx��
G��y�$�U4���1�����j���8�FYd�$�\f�[�Ї�L�2���A �ʿ�D�Z����+�!��,������#�é�A�\x�\���c9o�X�h(����(6�O)�)1�%�Ћ`@[7�߈M$sv�j� w�
f��QY���ml����p���KL�d�]�i����n���������L�
���92w�#�ǖ�?
Sf�i^��
Z���xC��rΈô�!n������%����l���:� ��x߳����:�i����D1Nu�q�Vi%G�}���F������|}u��ۃ�ƨ�>����hs*	����t]Ð�c<�3���_�ߞލ�C&���s�6e4|Ԇ�U���^�{r�|��W��ǖE�Ra���������	$&�D�;�������Z%R�8�u<āY�n�2E���V;���Z�6gٙ��M?Q���J��ur���k�M.$��qj��z��n��PK��v�Tf��BZ�V������fI�ۿ&���Һ����b��_�~<���CK�O�	a���Y�d��6���y:K�[���Q��޻&%�ɴ&wX<M�E_B�M�7l/(*���P�����1�b�!�1K�g%԰�`�C+���2��O�8����kv��x8�װ���5��01���&��G=�}8t#l�¢���v.�6'|��@z�E��#$��11O�rD�#x�O�RS��(5Ұ� }���4�p�˨���bQ8�,�M_��แ9��v?�WN~'�F�T�]R3�N&ѓXgnK�� "�H۰�w?��L�^v#ߦ�3��v o���N�X��>U�O�-T�׽4��ȕP"����L�뗩�v�Zmh1�	��h�����I�
���d����fziak�ա+�dV���fc7��S���T՘�LX��ǜn��=2��a��2���)��Ѫ�oj4�h/���'Md�A� �"���{��;�C�'�u�  ����<8�ow���[<��k���T��L���{s��vto�iA�D�¡���|��u���,%���PYc���m�^��v�b��[� 5A�_��u�^���	�L'��D��{X���9]1�N)���à/�Q�$NmP';b�|��5Aza'ү�rO�"�L�����J�� 5w��z�����Y��2�*a���t�:rMPS��*��V'�`\\�P�����e��������SPm���3�@��'$��"-�4����X�'5 ����&s����t���{�GՒ~L��m�h��K/�� �`)�� q�94��x�U|���^���x�ղOCeQt��R���њ_� ��1�)B1�*���-���4r"\H��]S�CG��+���Dd}T����hFY�p2��YqKg�	I���C��ZUA1QI����~�z�Jqi�����R�/�z�R�S�H�U��ZC�"x���:aX�8�I��G���d����f/ j�,�du!"7�����+��Rz�Qח����d�������8n���l���O�Ո{�44�_���Y�6Kjh�N�>kQE0]�2Vi�!Hإ�?[�����)�c�D?�٣�1��ޅ��I�B���2�0��b��O!�v\�$�?� ?� l���FP��PB��a��,���l��4F�ns������)a�;�Rt��p��Pq����� e�S�#��N��W������a�ws|�o��Oq�>�M�2EacXMk2�uъL�>�H��v��B'����s��ڽZD!����@�a���X:Y0�lo_�p7D���ߗvݚ�.h�>�P�)hv7���6X_zM��'f,k�2y�c������/�OS�ҿ�y�� ;�ٟ� `�� (��gs�&�Z�y��s]y��g�ں'����fLf� �c6Gފ[}4���!���zn����<ł��V�@M;E|ϙ�~�OLi�DUY{\�u�K������&��hs�J�����J� i�*_Yn;�*�3�iy���r�(��O�(u
���ͣ��(/V����)g���*O��G�e?{#%��ԣ!��x��x�k�\.����@֯g�&k������mH�q;���+�Mi6�%ww����oc@�4�� ��ɪsA=�;��M�����1���� �x㯣#�_�R����7�%��-�P�;��Y���G������ݖ�a�:k�M�s���\��3Ʈ��ۍ'�@':�/'����b����%R�M��"8)L�Ma�[�d�~u��`���Ƃ�&��.H'����H���Fk��&��~Ȓ�o�%�K�<68����J��p�w���.��^��E] ��J՗�KȠSQf$�5�9����<b�X0;�M!���k�����q^A�����<�.��ei��n��b��{;bC)�h�i���a<�I�7�6I�,�������^�SZ/��;�S�}4���BY�i�Ԫ��s��Z��@D��`����܉�����M�_�y����6���[����X��N�1E+|4xz(�]a>�ͦ��\8������{�"do�\����%��U-Mp�������rf��!b�.����b�q�-$�oA����&���Ѽ��Fz������*��(ت��W��]>y�?$����	�"î2]��I���
x��w��.) �{^��Ѧ�ɳ�rà�룴S�w��T��m܍E��2�E�١��\F���c	���)��2�r�I�J΢3}�e'4(dvDK�IZk��5����3R	P������ѹ�1ƪ�@��nQ\��^+?f�a��@-�dm���Ň֑{�x��ɍK�k�V��("�׺t�ߵӞ�]��CZ>�:� ���*�?�p=�������L�4����`�&�o���k���!H��ӝ[��]n�_C��^/\&ܻ`�u��ӿ-{P��3w���#��
�QF�w�
lM��04I9Sja��K%
�i�6D&X�j��nzQ�,/8��R�r��Ș�0����{�I�����v�X� ��0q���q�gd'���)Ig����%�S*��,���@��Жw���]qd���v��p�o��|��0�j3��-������^ |��]h�ƥBt������J�%"KYy�ׄg1nɺr�?�O��T�uЦy.�e���_xw��#��u΋2E�C53O5Ǫ�p`�L�U.s2�m��wI4@y���E{3U�å�QO�W�y�h'�P۞���x�G��ﵐ�s�
j��>���-��3v�󫀌�^�H;��3����w��ﱑA\ և�CV���PJ^ʉ��dR�R*��7� �xʀ強�D�����Q0#��a�ʴ� �вכә	��,���fOj��Cҳ @[������3�ŸYx
u�4�r��Q%v�z�)�
�\�5`��,�mQ�!Đ�����g��X�4|[+�/�q�f�f�@���*)!�Ҟ��7T����p�����{�&;����Ld��5�W��0E���@���� �^�A�Vw�V.�� 0y��?��8�����9X�<K1��W�#����"��,��	�y̍I=�k�Ha�L�gd6�]�D��6�lD��\��1~�݅D���b�\�%hD������|���bwB̟�U�u���<�UΦ|�%H�^��V��P!:��>*�����Q�t�����J��T��3ݶ�gW��0�m+����[AVo�ʞ��/=#vv�����%����>��3���?Ψ��vC��%7��oڮ�XRyW��=p	_�|��a@����L�EDŏ��8�)x�$�DN)�
�'�w3s3y���-���c����(��\�r����3�i�DP��P��踌�m�E!�0!�~�ti���Uۉ�RJ#�N��a1o��-��/c*/Eaw�3��-P�����K'EY����{������Ά�*3�H�/���U �y'�J�G
�uǱ�[2i#�m�Y���~-�i���p���~�ˢ�g�Q��.X�e������,��b��lv���aZGNވ/0��1�#�NYy�`a���Y/��<cjri�ӈn�F�� Oݞ�<�(11͖h��)OSN�@:��{1:-6S'U��Gt��O�8�q�C6'�0(M-@���']\*� ����=f�A��t����C�x�C�d����G���^�G����k���M������������r/V����/��eW^��
�|.6>U҄G� ���L�Y��0�O��5 �3��� �L[7��OH�8�e`���|�C�\�ڶஅ۵���o}8�9�8=V7`�JL�|> C�]fPU6e=��pp��)�����f04�FG�s^��n�C	��h��0MrF��B�Je�W)����[���EW{4�e���]���{u.�5h�E��H��(=��;��a!��мdJo���9�l�j���m�d|:u�w�3�G�2nO�a|�7��8z,e��c�v�e�N� c�ei(ٻ�������Țg����
�����Y��V��O&�<˭��Ѿ���4�݂;:���R���#���i��%��,���J�&�z�OoY�[�o"\�v��S����P�0�h�;�ORsv7G]"�$�诺
�Q�-M��[��l�"֘����{Sa�}hM�C�ꎟr��M���F3i(�)���!9Nl�|�;6&�QH8J�7E�!��=v�-��J$�"�j���5��K$�F��.���W��?
�@��&=�>p��ͧ�ӚA�:�"+A~�4�������iz�^�[��o!��y�۰T&�&\X��	��������q��Z��"���h5�C���Or��r��h�e���wq�Ⱦ8
E]}��!O?��
0c�;'�=ƟS+|��:�Ε�I�i6V:���ۯ(�T�J���ԫd���L�l�f�T ���|�GT��-u�����W���u8Q@�!l���}�����TF C���NNET��\���|C��"���k>4K��hA~��}z���AgW�㮣%�#����+�l��H���V��QP��I�4��݉٫aP*b΅Z����C֍��
Ěհ�Sʲ�-&��.�[1��P�TBl� �sGS_��-=�#7���L�@�`l^�Q
D�8Kʺ|B[�,�	���w%E)n[���Kj��C`��c'{b��OB'���[*���QK�kl̈�M&��J����hyG0U���!ǕU�ɰ
�I���{�ǥ �EpD�"������l#أs����AvTbo-�q���ݜ���q�.���м �L�@m5u�<]�K���UV��/7������B�y �h���k�TȄ���k�٨ɋ�a���rֲЩ�5]}��vw
2.��t�U�uJ���(H>��Vc25������\�+�n{��:���XoB��fR�2�v� \D��$�`�<���o�=������ͫdx��W�ljڟ�,�+��A����ޛ�֔��J n��Ңd�0y�dL��Pf,؈FȠ�e&&l��I��ȭ���M{���&�+�o?�R��e���`��{��E���	�ոE�ɴ8*E�b%w���^*F<�տ'i��}f�$�<S��v�۠\�4�{?}�O��b�AV�XY��6�_p�Tdb1
|&�L���m���e#'V�w���[�X��8��l������p�_����f�d���"��؄7RS�j�Nx3M�����v9y�Ƕ85��e@������ზ� ����P���Lf�_#yF�h_(�ħW-��u4����;�=X��3v��~�بY'���@��6����0ePW��d�`QG�kM���\�#��]���߿E?�^�$=���+���l�[H�)Fq`�R��sT�u����LBtb�KjI�|u���D7�z��Y�)�J�ʔ�!�!������z���}�C�<3p�LNNJ`��1z�^�-ʏZ��G�}�/��C���rG�=Gf����:H�˩��i��%��m�-^�䐎hə�q��o�I�ZHa҅/�Ї���!�FS':�A�' ����l��=�0��W���a� Y�3�sƍ�m2�ix�/n��uA�9/0��9������*���]���@1��0;��\���-`	%5�� �.ŨR#��pW{�dJ@��a��f���);@͑�w}4C%a8E^f���U��O� �|��� �/@����յaؿ"���mf�󮢇yb��ܞ+�l��
�xm&(�얙e�#Q��F5U5>?ǿ�y���OMϊ�z揇��,���b>�c�;琇�y9����q��ت!�:���,�#�|O%j@MX֑��8}��w6����{��2ެy���O\k8�1P��7���6n"�Xe�?2aF��2c��!��PT9)e�)6%�b��A/3�����u�j�ɯ��D����S�p�1:,�#���t�*���x�+���F�������������-�ZX����^�En���i�����P���HQf�JG�Ҧf�N� s:��#��x�!�0���Բ�F+	�l������ݜ�������#+�m}�(�N8�*6\pT������(7�^#�x9�~�PX
�L�q����"�RF�.�6J�U�(O�����?x5�H��Z�m�a�����5��Mř�t���@i��c�4�=۪�F� �P�n��7�l�t`�g07n�f��P`I�	s��{��������dB�F��p#�ł�4����}��S*f!7��踹)��m�䍰A�S�����C�v�W�EE��j+ ����XQS��;��V���Mb8�@Uy�罗���\�5�̣R[o����$FI˱󟲦(�\JÒ���{���h�[S�+M2�قK�M��J켛��'�.�\��4a�3Bn�>9�;���>auï"1�n�C0��($R,3+���
(�N��CU���]�����*D^A��0�)��kTF�u������~h�VnB-8	_��$�� �5�v)��d�����ЕY��2}�p������>r�u��zg� �h1��]��_K4�Baw�����3h��߱� +���m/��1�&������j�5��#]����˧��$�h=�^��ݯ��Ǵ���i�@��,,9r����v�)�P��;�s'O��L�b��$U`G�ǅ�ϖ�C�[Vf�3��(Q���Y5��s���P�OJ�:�:G�����0�l���Rʩ[����]�#�7�< P4Nє�A〄��o>��m���G�������^��<wT�	��84�I�~8�9x�U��[�畯y�O��S��%�gH+5�&J''�����bi��lɼjJ�>PGУ�-�Kzv7ʕ@^�YҎ�)Zĥ���9kd�~cF14��^4�� �T�~�7�˟���2���7��pqT>��N�p�]Ʈ��=�O����'�V@Nf��>+/���Ξ��B����z@�6[�ˆ�<xh7I+��O[�06ޞ���\p�Vv�|Q���Ƣa����l����ץ�f��� ,�lg���I 3mg}��(5;^�~��?�:���ڽ�O��+'��^�P�y������u2"b��%8������ž/�������QX�c7�>�X,ö���ϫ	�iiy�S�a��J�K�r��ިV!��)P�$�H͌�n�>�]�#y�菸��<�ⷰڠ D��醦��Y�">�+;��)['¤�eh5ū9
���$,�C�{�J�Ke�5��;g�N��JN_�ټ�V\�K��6��7}%q|Y@u�P��-.�F
5�`���s���V�U�Ȧ�����m�Q$;O�׎o���٬��-�yX�8��ؖ������w�ͪǸ���D�ؚ�w�g�� `4�,z�b�nw{�i��7#Wf���$�_�=��Ը�lY�#�3�
G�J&/�<G��T�WZ_�K7'@�]p�,��1Y$,-\�x1k�nCm����`0�R"G>!��#��J��ס�����^qk��5~�Q���#��`�UmPTB�_�)��l�5��O2x��a<e�S.�,�a�&V����Ģr		�ʷ܊6�7H�h��tp��R ���B�a����!E'l%�ع`O�5?� ���S�&1�z�0���y3�mol�c�2<ˈ����t�OAa,J9fᔏ����2�߃�Lqf�Fy��!���|�|:��Q,1s��#=X��~dƨP��������p�!>Tz�� a#t�рh|3�>8o,j >/5�����:ܼW�`��6���u�y�m>u�W{>��J�����;J!���9��?��0�Ƙ�o B����ҿ:�H��5�u��!g�uL*��H�+�h�t�:v�u���2bR���QS�������ǾI�$?�������y����F��X�������m֜V������|5�T��1s?����Nt��U�j�z�'����^lfzjcR�i����}��(N����F7�6\!5blx5X;��^�~��K�ɵ�^^W��-�zNI�7��H�U~�^��t8#���iįG�ȣE�����DE����=��I����y(�dK����k�v���ȭ-Vd�ZLZ�~�
6/�ap(������h/�� Pa1n&U-(�p�C�������z1iKj�⪈�������Au�Vm9q��r#�w�g�Āp�UHO��,���7)����)�/�������UZ1ѵ(u*�U�.�n.����1~0{�w
Wg�D�ZڵR�G(U�͐����R�D�X8�e/#z� �⸍)�X�^us�����J^��l�7N-��c>~
P��:�d-����V/����/]��C �A�����םߏ*�s={+I�_mWKf->u� x�w ߂A��47/l��%��+=�?Z��ص�6����JIc��� �m2�c�H������I�J,�*S{+�W&���pGxǒP��,�,-�[�(��,U��*����v���Bw�ъ��9�h���[D���z�_�;���.w�o�F	f7��f|����8`��,���	p1��i��{����Z ����g��������>�|��cS ��T�ʚ�hE�oyukC�}\	k?��)��-��r�.ލ��|]�ɭ ]$��IU�aB[*㾵ȳ��x�,G���"�j���$S}��'������]����Jw��S/�!-��8ێ�-{���exiU��a�T���1���4�=�=߇<�Y:����[9榓����y6���:�G4�	��Ru���GM-��B�9�$]��4��)�[Y����~hϩv�d���t��f[�\�^�=Wִ�cl6I�pDk��A�A��:,�q��M��ö-�r�\��H����)���B��`ݳ�(z��͙V"\�.6W��S�J��lԀ�.��&�n�h<��'���a$��\5�������8�g������¶��lc�L�{y<�6]�d��d�h�|���bM�*	���)�:5�h��۪N@o�)EL������.\%]C0r]�/��7��`(�58¢#lڸRhj<@�R2� �S7T�X�Yg~7�2��\���v����zSJ�؞���ru���V���Ou��֌�q�o�Ѡ<Y�t�/Z3��t`���Ӊ` n��F߸��te��*� J&:�����+����:R��?-�h�����T����D{����;��&��3]1�rr5[��Am ��w�������������Ϣ]z���=S·�&�𤞰~�릋?��b_$W�1�KkI[^]K2�mvaPr�j@#��ڦګڃ�A��{͜O|�)�"�����"���jk]�v���Ӆ@��PA�M��,A��(�b`�5︜����
��0EV�x�Z/�F^*'�=sبr�G%�)��m]{Z�׊�\��Ch��ZC���A<�|~&Ǵ:">6+���D�i��J�h=UŸ8ja� ���Q�/FX,��C5s�����ܧ���U�^X��;���ca��
d8@�yi�H� �9B��)L<W�(�.�i��������q��ەr_��݅��t���{�dZr���uD��j,�k0�'� w�j�᷈��af����~�!���~-�C�_��m;���r��k��֞���_���Va������Fן� ǃ�����3H�����r2�F��@sI&�Fi���:"�3�H�	J݉���p����F.��m���L�E�
��{'>�����;�z$�l�xLU������Z��x"��߳׈���߀��c�cl��яH ]?B.q�%����J~W�<��~����6�=m2�Ci�U�ܱ��5��m=��In#�w��������9b��湄@fކ׋
6MI���]KG�3��Q��̬[������v�)=��������sHֵ�.�d�����ңqn��e���G���@,٬�s�I֭h�#��Qq�/v[��[�QI{��U��J9
^���t�Gg�+^��!�Kr�&fj�J\�%4���/���7�``�v�(���O��]|��N	c����h�T�P+�z-ǋydP�ش��\1n?�P�� ��Xq0Xa�X�����)�&VTbb��3��<�[z��Rƫ��/Eo,T�y�G�Uq��M���H��u�5���:xN�l-��3�����Y`PŀF^�Z3H���}kX�#)| t��?[�a5��M*�R��R�X�|�7�A��W�$.���7 ����
�@vJ��a�	5e}�B���'�T�P�i#�1e�T�z19�����7β��j)s��Ml;�<�T���-�?��� �~u<�oi���X�袦�ڻ��L���-��焥&�o���p�݁���S	�Ǟ�Ǝ35d8�	��p��o1Z���?��	�<\Q��k����������B6���)3���ÈO�F"ޞɢ����s@�����_�-�1j,<̢��GU��wy 13��x�?��2I�k4�S�׾	K՚f���0x3;[��4!%)�����L��crwy���ϧA�<QHU�9�D�4{hz�5 '̭��!� y/��fY� J��;nP��-��q����x�QW�>�h)c9�b�A:-����D����.�NT��ѻ"O�]ȁ��pd_�=��J�_k���^�__Z���9��#b���δ���6@��o�(��٥�g����y�%y؅�x'!��|�yb*o�N�(Ȝ"���*��9ѕ���[m�q�[u�.F��~��>3�#s�j��T`'���i;tTwo4�� |�)dFs��Տ,�/�PU�f�q@���ك�$>t�V�意���]�Xp����'��s D����.�?�S �1$<��<`��͇p��k�˅��fd�z ��nێ��̹�~Iߖ~'ҹD��=%)m�95�tJS�rضl�  �A��>�A�ٷIn�z��1���n�s�a��4*��r�߁Sf9�O����a�i6BG��JJ����/�̵� u4��I��vQ+�H��a�~�b��W�@Ett�JhM��O/� �9
�-��
O�}�93uu/'`���qQK�A&�ĺqR�xa��zv`eA����t߯7H�n��2��|��;����o�+�(��'�,��
	 ������6�+`Q�^����Cm���Y��9m�ܽ��A���7�g����8�gp;f�)��RZ-�I�א�p������CG=�J�^s} �����9+\��O�{�9(�u:�^e5�#��ǐ�}+2Ga�u&Y�K��A˿ص�V6vhR���)c��ΕR&$8o�ԧ������s�!h�s��Gr�'����լ۟uT��uQԧ���BF�JBnxl�hAO�ufģ�,�&G=��|j���j���,��f{�Nɟs͒e�J�a�ğ2W*s��Q�3�t�i�8O�"�APzXvq�.������X%Wa(y�XȪ*V�v���A�7Ezf@xpJ
�`r-$��� �l!|��W�c��36�cyh"�N���@������)��Z�!��WD�B���1��,�EK��(G���3�9�ɀbg%��ZL�*�o���޼�iL���Hfl ]�e�6 ��n�-�r'�����}�9U�`��o[?E)%b9�s�g�%���hߒ�)�֛�5Yo��J� �d�C��R"��l���iʦY@����Hǯ��
��.uşM�"�� ��4>��	��8ߌ����Daq�&�+cY��9�3�b�|.�F�n�^��I����T�Xþ�ᇝ�
ב%��&=���K�ߠ.2ɰ�/̝�\���n׆6��"�ҩP�ahv�f�1"B���9�� P\�����ϭ���X�=o���%U�%�o�(uLN8�z=��{�ӻ��ڙRb�����J�� �l��w`7�9�|vZ�B�A�K&_u�)���?L��(x>9����C��)_��jM�/�FZ�����'V^��1�j�%��轗��ű?�r�`�#�8ׂ"NE��Oe�-d��.̕�Ns�ڇ�Z�|��֘���OƻyJ_$u�><���t��®���W4J�k^H<�Wo1��]��v�K�a�a4,� ^[е�<�ٵ������$���)�SE���)�T�%a�nHK�Lv�Υ����l|��������MȢ��C�*��$���e�$y��=M��g�W��Sd�����hL/�PF ؜�������pڑC�M�Y���9�3`iJ�`L����#}��im�3�[Ww�b���.���r�B$`���T��
Ѭ���@�*Ҫ�Y*��V�{�&�E��B#n�X�ʬ� f�q��t���vw�%6	z� ��M�rGlف�����ʸ��Ӎ��sFhE�M���e��#\�{kF���O���(�
�)����&�F��Z�[b�5a��&�-e��\��o�D����C�<u�-,[�W�x?"dn\�z�����EKAEJCQ��9�V�z*t����(�ғ3@|��`�|�[� S�A��v0Jd�J��@W�ń�>�Q<�{��#��!W��m�ҭ�|�$7Dh� ���0W�4;�y=k�(�=rqJHVM���%"]�!cyy�W����TW���%�؝`O��o���]"�ۃ8E
��?���#�E��咩 	w,��U��Ш��m���y�R�o��%k�刯�@>P�߫��g�7�����I��I./npܱ0n��Cu�*уnfF��tYX��[pĎ@��V�ց6,t��v%utR�-������ۯ��܄�RaEr�݄Q*,�X�Ǒ��ʁX��y�.lj���m �c4y�d�g )�o�ȺF�|�|�f���@������S-%.&�c�t�X�Q��~�m�7}�q ٗ��b�!s!l���" W�f���ɽ�c�c����>����]�^�i����`�W��	i�����_>Ώ�ZY�?�Z�:}"&A��̡�l���צ�\OH�P�l�+z��}Us��f�iJ��W���БP�ꠘ���Ml܇\�' ~�F�J�T-����AȩB��|��7|�df�iR�28��\�7�������B��l�Chi�v�ہ�Wux0ᔖ��z�8�R�!�t��D?�PO;�xچ?
\��lmoVՙ1ب�o|:^������[Ea#2��an�j��� �����p��Mi�����d�]>�����k����QY}�I��v�τa�,,�8-��U'kA����>y&�����>)��F,<E�X��x��Ռ�Y���է��A~��cl��@��>⌠ȇmłw��,d�KR4���A�W�:�h0ϱ���S�o�e~�ǩ|G�P�XAo� x:&*���䳷������S��$�}ѥ[�ֲ���}���EN+b�����������)p���_�&*�q2
{B��C3{u��<�"8v����_������TT��t���V��Uvïja_�6��U-��<�"���LI� ��o�C��l�W�Y�0���2���3=�5H�+|ִd�ic�F+��J�p�/Փ��We���������j����_���IjxIeЀ��>3tı�L璘͊���Y�Q�K@�k�ѝ/�Da~�&��L�?�C�G^@$����Hy�	��O*��I��{������F�[���ZKfJnqi���Euk�^vIFet'����b��Ž�R��ND��a�ZK��o�}�:�sqܝ��m��to��`18���#�A�P
�$T��x��.���m������u����X�4o��$��%C����K:s"�0�4���+i�b�	��,}� ���n"A�
1�R\��2�Ė�x�%�7�&-��4���+rFq:s�ϰk�q�Ne�<����A�z9��2{oeANoj��3���h�t!9�./�'p9���ޘ�i���A����`��?9�.8l��D3��C�����ڗ랈ŏE�"�"9�+�0�<D���!�y��W2ǽ)��Y	�l�&�o�iQ�e:��Ď��P��x�z�jD�0�)(v���6if�i�Ea�M M_��#\�ON�q|,��,z'�8F�=T�xbK�I]�P��[[!l"�_AO�}�*�a�hgJޚz~��_������GW�޺�4�@�'�_u}dwF麁 ��=t��ډ6B�8����4:����g!m^��皖�蜳�ǂKxؕ���� T�a��#�!_1%��������^4��5H�7p��ys��qD��O��)����7�L�źX��sp�)�梙��(@2(�(�^�N��K�	�p���s۰�D�4��E�?�|liee4���|���ՔCN#;q�ckn�s��Kه�L<�N�'5x��=���ܻ$�2�V��U����s� �l�{_�l*&xX� :UD�
�?rCM�8��[�yΨc0����3���\ʅ��Z'�]���Rv�Y}���xC�kc��+?4�T��]oLe��Y�%<�ez��Cn���|7{�qPE��$RǮ�A��u=��5�(�=j���tƪ����|�ML�o���0�-{���A������E��/��X��-o�ZF��X�d�F�&��v�Rє1M�ڎC>\��ok�;��I�j�qOD�h&��6��!no�F΃J.�oԇ� ����wl�x��ǂȯ��!�O1�t�έs�_g�@�HدѸ�� ��.���s�eaѕ���v�EZÖۆ+F+���8x�ٹ�$�ehl�v�ٴ�{k9�vC�Ce<��zH�� �f����v,#�a��?il�	ا�@����rО����!S���r���F�\ �C��u���B'� �i7r�cK,�J}p=�d��ˉ��2�G;��:�[�-��M�J4Q@�4���"�&�|�g�H_��v)cF^��M��a	�����vnZ����y�h?��T[��%gK��;!�l^��㧛�	�:�SF�l<	�e�4�j�0���#ES�[����vC8���E[��e�էa�X\NF���I ��®!�^!q�T���Y�U�<�s�* �rs��7���/��bz���:� ��qq��}� ���6-���E~�"�&>��3V�����n�U!_7�I��F� �yi���@���9�Q;E�������������{����g�X��� m���N�[?;{@��u�2F}��i��#%9��N�ВEr;PO(�%��K��}n�Ӝ�A����F�D�7�����
�t��g� �*�!��/ud�(������ᶺ8�gz�����0�h���t��&m��~12��抶h�.h���J��<�y
���F�2����ppIJ��Z�u�V����s���y��B��D���k�.>���+n�w?ۗ��m���v��%��Z"��V�~=3��#�K��y�_����D��ɏ��p�Iw���G�&*-��p�:G��ht;���7���&��\5X[������s��F�n<�W��i���9�47�+
Ce��r�>���}�{�PHcX|G����a:e��B�f:��$s�E��q]r�P ��ؘB!T�W�����M�S��ݣ��*�k��Eǅ�A����Y!�4�%��E{ޟ@��*U��A��ceY6���5;A:O��k��nz
�S9Q|C�ڍ9����@ךY�r�S�Ԏp�B���}��P�|�>�^�@�HH���;U���:��/�\���HJr����l�q��^�oYs�Q�z��<�f�v��wDwp$�(�<��_��Q����q$�̎���G���� �n��t��o���G�5��T�P���S�~8T���N�:ߊ� �f�猐�+6x��n����ۺ�`#���lz�U5�,u��P $ωm^�VymQ�"r5rO��)}��O��I�t�v/ۛ��	�@zH���H|Tō�λ�9���hm���qyX!� +7K�!���șt�� _D����u8l;(D^.�И齄tg�I�a��H;x h0�N;�AĴ/�-��`>�jF[�&7��'5��D�;�:sf:��Oi���>5s�{�Ţ����x ��Z����4f\}�>�u��O���Tɹx���R�kPok�F5�Ѝew����k.a���V/�����<b������H�O�8pX�=S���x}�}q��*D'�p�}��=����O���.1-Q0�:Y$���v?B4��2G ��cr�z�SM����H���t��<�Y�xk��H��Fm�p��EK9ĉ�M5m�����\�W�\��-�4�?ߪҶ~� �{�B�PI�a�G�T�I!���Q��ѫ?B@>�GOE�M��{�h�Q n�+�v�| jD�S�
D:MЫ�;i��[豍�\{��k :r���iE1�8Q<��[A��ح�0>��*&��j���$����w�P��<��9|��$�?=.dR(�����>����Z������]��w�ivq��APP�C�rIr�������p�"���@�Vi�D�)�#����v6zxWk�àٱJ�}�a���JK��s�ۓg�+��ɓ�w�¡\"�T��}��������-�`e��ʦ�&$��U����Z�t����Qm�t"��f�SB3�	�����Š�-����	���J�1���|���[w44�?\�%�4�2����T_�Jj2`�)>o ��0g��a�L��få-)4V5��X!pe-V�W��~������r�3�zOd�6���?�bV暈^�Nś��R"I8<H����)�c�)ݥ)W�����6t�#���0�zV.��5��'6�oIA����ɘ7�6�a.���ȧm0���({)uYA�c��3��b`�u.�YY�ߑ�F|�]��.��'���7�+��0���<z�P\��)I��H��W��W��ŉ�:e�6�t5�a����A�U���Y部�GM��������Nߢ��u����ȡy5�J�d��͔�Y�GX��p-8��arg�*���oC�9����O4��~�O�Ȃ4ΒA�=l�2U� W
�r%����HHj����9�PK��vA#R@�	�H�
���Q�*ˌ�1Z^$�EC���h!n!E�X��;�wR��j�(�t>M�9�)!�Ԫ�`�0(yk~Ӯ.k
�,f�/���JN��Wav��9��r{I��}%3klb�P����=��{׵�+���PM|X�������l�ТށM����\�� lyr���v ����m�Z��M�����./��Wc5�Ŭ�W^{�y6���\!3�śk��OB�w͊����</�}�I҆	U��0;�4�;p'W�e������0�^ Ԣ�񏌐�s�`μ��{�E��X��� ��,᭙ۄ���3�U�h���37�s���PB޽�����!5}S����*v�GȌT�C����oN��kZ�"w!�2���0[~���N0?@j�7C"����`:�ч^c)��;|7�ق|i3�����*�t/��U�
�GdU���E��0ֻ�����d�a���̪Fb���A�Ww���5��Ϻ�.&�)ߍc�kG�8-����h��d��%*JXJ���(�X��/4[;?���L�_G
|�8��u���]�K���o�-��M*�S�4�$�}"���W!3&����A��ܜj�7��Qez('��%��䟚����*7�~ׂ���3�<5C��X�gOj�?��Yd�.1�C �>���p��΀�*l���sXW�i�q 2)���Z�c���;��PE|"I�1�Ȇ!�I`�f>H:�*aE�uD���_��'��hh��j�\ؓ{J@O�����.vQB;��3�<���?O3��EM�,�Ѓ�U�1�P��;bf�=ȭ?8��y����退{)���oGIv�L���:=�9�A��-�m+@���ӎL	)	�Xh$��#$�z$��ژ���I6�5����L�L�L�n�:[��2�����AB��c�a
����SJ�}8ő^��ǣ%�y���696���j����ɤ�И.*�R�Ib2��q��Jt�x
Iado�!���}n����
��G'aɥ!�FIʭ���0��{؛?�l�JΉK{���#&�@�'-�@*�^ ����"��1`���{7�C$�{��<�Ud ��g�<��?珓�"��xl4%?,NA�G�}��	y��f{}n�T�?;�P
�{H���2�]'�vR�ƺ1Z�c�Bɯ�Dﮇ'�h�����XH��=��V�rM�8Y������̅�K)�|f�����]�J  KJ*^��Sy��c���Oҵ�T���Ԃ
�V�LXn��*m$c7\ؖul}���������@��6���n u~���f���=te�d"��K/E���y�T{�)��t�b("+~�vU*W��.�BP��n�ңi�MMdn��X�F�>��הx�x��۔�
�q�@I��"ڟ�m�[��E6AOEI������fbk�)��R��o�*�Q�j�� F���|Ow?������9LZ~R<C$S���i3낛먡�$:{��|��Y�ե�� s8�tq�M!�k�F�A���K��t�o�/�	���j]2{��0���Bcy`ڝ��Cù.��X��u�hszE������j��n���y���(&�p��*�X����;�qx�"�yfp(+�n�D���V-Z�:i�zq��J�o��N��O��b�p}�3!�y,��39�����5�o�����&/nzd�J��(0����;��Z^ݍ�#-h��"����C���L?��=_�����{!�>g�p7��X�2ʠ�'��l��I�r)j;Hyt��*83�v�����Qd���ƛ�koSjH�Y�� ��֨>P̷�<:����<���N*Ӥ���+�Xet�%�z������g�|�"��U���}ͱ˜	��0�@�b�Sn؃$
q�ZM�}�&���=����$t��9^d1�j��������-MuN��d��]hL�=��y�T˗�/U6�2�q���B������B�4\�q9I�6�����;Ĭ>3o!acS:�%�<98���ی>�.�OW���Z�|� ��������,ˆ6ʎ@!�5���π/�7�RbB�y
�\�Ѫ�~�3�}��g�""�J�U�n	+��;<���%s��ٮ��S%~�_�3��1�̄�v|�p�\i@3'#O�_��������9�Zerݖ�������*�U~���_�n6qǔ��*w����y���D+#;�}u֨Mlo�M��U�P�ԯ��\53E����RX� �R�id��Q��No$�:*9��Uw�?�k�@D��� 	����.W��6��\;?#C�9�_oE����3�炌��T��I�B3���S��+���ee�֐���G�h�W;}�K�=ZA=x۴��͛�63b�8�)8�N)J3���&����������90�W�/}*� ��i�w��RJ��*�c�_vY�=�:3G
��ߊc��+gyҔ�/�(#ta����-��t*3�ii u�wx��j�],�u2%ĥ����Y3�܀/_��hUN}4�`D� �8�O�du�jAL"�1G�K�CF�QB׋֌��4H���gۦ�2�d:�s o�;��M	�T(����S�:�@�w�AW8m[ve�5h)��s"���7��$�����2��u���m�Q�,��=Ɇ~���,��.� c5���2�u�|���:�����i���x����!�M��U�����y3ԈX5�`���7S9uDH�3Q1]~�������p'\j�3��w����~���Q|��A�n��ϫ�:���֎�e�b+���zc�BC�6�����`�HG_Ɏ�nc��+zQʵ�B�7���l�+����A��N[T�@��e��8��'_M&��{�>s�TG�����Y�gOH��<��@s��	lZ��Ҥj��utk�ɽ'����Upb�)W�dL1Jz4%���ئ�}�٫��@�K�b~��%����U�nx�v@�YW]����)P�)-��f�{f�'��*c�,=d|$�t}!���@�ad5�����ώ��;K��N
x��d����R���{��� ��f���଑�
�O�Ž�,M&[F��m6�/��N�rWX������������qGȾ[�y���m�~���Zd���HL0�Z���۞�qȚ�m�y}�>���JΕ�롅t���u�ެ���������ԟ��E�S����>d���;U��g�%u�u��g͌�R�n�:!���y�|���x����I�V���m�7�]߹)����V$�`�.K\ ��`	:,[�I��L�����g��a��5��^f7+����Y���s�*U�ѵȘ�R♿�d�{�����J�;��5�%f��GB��3��/�B�,1�y�kH��Rq��S��^�`���s{�zdZ����d��1���p�ɨ���(s�Hj�pUY��&�/��[�_�fK��e�ƿ6�?��:���@��ӝ��D-4�ㇻ�V��&��}Z7�"kq�'���`�w�̎i�z��U�I��$�����2M��~�uZ�p��=uk�Ub�����X�,D��������>��a�U ��@�Y42�ŕt������\��2^HXS��f{f2����8ߡ���%l%�tQ�O���X��j�_��� ����U� ^~��.��-^Y�ZF �>*�`��>�y�����J�m����R�X�h?s:Ӧ0��ں6
)����x���\��Y H^���[)�<~�3my�J�1'lK�U$�g��c2�3�lR(������*�>S��)����DQ�I]A�`]���a�#��/`x�qu�sk�� ������]D� �I���Hr��dT�j���6)������D"������]2�XsTG���9d+�Ө� ����QU(���C	�9�� �%xaS�E�vISB�	�AX�_��mG�%�Ѻ�T����^x�<���0�� �������A���u�H(�5F�ZߢiKU�(\���'&~2���H3�>t?ȡ�LbB򪕐T`��r���O�pt��s%��{��-��,ûm��qp��A�ۆ
A�d��w6?��d�IW63��@��h��	[���O	֧���/�tp�4��2M��Lf�Ð���Z&�����+{�b�<�i�!�u2%��_��>��T�I�7M��>�e�*i�"�]!vu�<��
r��B&)CA��gpa�
YZ�ظ�ՙ��e1�X
��c��^��Y�^,���{/���4�0�e�b�Kr_�c1�T�\�@;PAZFNWJS��Ӫ�)p�a���{ނ<k՘�G��13�=�������k��O����^�3!ΐ�K�C��4���M�1�}�?�($��"hT��̖H� sW�=E�KkeC���z�A ����[G�&ۆ��[-����zfƘ��)5f�����
b�|��U��v;g�H��Y��}eùk`$Y(��8q7��8��>�͎�h)?k������cXgX�d��E�FEt��D T۴>�����H5�"�?�X�.'Sj�<G(���d��m���"U��I��&��Y������	�2y��O����gt`�	��܋��ik�6�5��jW!��K� l���L<hXH<���\)��P�1�N��B�(�q{�]4��O}�Gv�"�j�'�s�T���0XWu�8��U�&n�;mfpj/Q�MÞ�]81T?f���l�{rw��Xv8��<�i��������sr���9~�>c%�ic+����v�ޔ�i�d�ox�mk����r~p҂2+w�ͰN�V��ܸ��K���[H�W��1W>X'�c���P-:cSf�"V��q�&9,�[[���Bd���23$b.��W��5��<}⊥U��P/��0t�oυ�%���lf���|�N5��$w]<.�ZZ��~Z�Q��N��ATgë��C�b��w¸�cP<�'��}�3���s\�	�b��K�uP�2p��F�5�����M�����6�
�}���BO�������GUn���J�Ղf­����?O+5���)R9�9D"�4 ���A;���h�ж���T�C�VH��F�2�}d���)S��G�)�Z�Q�*�_�	��TM"����\P�kJf���9#��ma9����Qr�a� _z�.��Y�MV6����f\+n�a^Y=��rR�D^Q�a�� ��O	�4���u<���@���;%'��Z�a�6L�s�e���t��ؠ�h?�����h�6�cp�Z.:&�$��@&�=�y1tNr�W^�d�ټ����y�Z9a�Rr�sK�d�ZXw=E�i�,��	n��*�Lsp4
��K0�	�u�5�8��1�єa�nX���ʥ�n���>2�u���V�R����u%����w�ƪ�LQ^ nj�h���s	c	Ob��(Q�|� ��j`��:Сy��X �K�/A���)��^��6���C�~~�6�r9(2yLm3.��/�D{<���嘧T�𔤬�-�N�F��.�c����l��b��q��C��/�j'�gM�5���t��fW���p���@l�}l狴h�' ���ښ��͍(N�>��{�����z�I�`�cf���	8YJM��-�\��Q$�Z�w>Aпb��	Ӥ
p��y�L/{�ֽD��ơI��5<���PU�!]��6[�2 �{������xW���y|����{D�z��EX���ؒ�GG+)%2ᾫ4��lB�/�K���}8���!܊�����J4s��1V���F P����`��"×s�P2
���FH�O�a�����O�Ue�lvM/�f�'�[�����Y���B  lz6�N|�)˦E,9��'�u��C����A;�������;���ӎ���i���{�.|���u�&�DY�l`l��'o�ZUZ_jT���~�y������V�fB;���-�[3	=�T��Nw�2C3a���rM�V�s�>m&�I�1/c %Kr Rk�h���!����=�oK�5�Cv� ��M��^��w�3�u@;#"�i�?~�P�j�:��숽W����\�#F)��O�/�	��:7�p��]�;|�R����J/�f�nJ��E�?�ʷ�E�VζgH�I��}���	F89r��Ic���{<���O��Z�)"�LkzD�� ��� Ź��B�� ��!������#x�ˍ���HE)N��N-7i��胚4n~L'��D4������M���X��L��^	͢G�J)|�&u���`�|�)/&��r��ߑ������ӓ���+� 13�t#�N�f8c!R\�c�:O�	�l8��y�&ǭ��������Ӊ�L#k����&U1!�ʟ����Rݓ(���s����8�g�q�&��#��������lN`��{�c9���5��T����E��MXv����pn%.��;�nz�۷�][�l)&�Ԏ.��Qʻ�QkՖZ�FI�����sPҜu��S�m㵣O�w�?Q�w9�rrȒZ<{�e�B��tՕwL�X0<�{�ͱ܍�(��.u�����2��.F�b��>#���+ �{K���5�F�I���)>��b�^��,�]��Q�-{��r0̝�- ��%����Ĩ��w�{)�� U�'����"��/hV{��
�B,#��g��.���k&n��55R���8�23�r�����u&��K#$+v�x�Xnr����>��55NJ٥�����I(��ȋ����u?ȏޢBd����Q�V��D��e���d��d��'`���ã�#+6�N�V���.����2�Yl/.�jf.Y鏯^m���]J�Aa���pX[r��拺�̎G�@)��WENq�s*����W�^�f�׭u05C�rq��?�j��
��m��nN�7�ԏ�g����Wlel�9ˑ���&@��� �s?Ƹ&d���R�|9k(���!����+����Gc+�<� ��'��8�5�k!�J��C�V��{�@{�1�=�d�! ��NTF�4�{����;*�iA��?�L!f��.�Z�ġp9�����%!�5R1����f��b.`lHM$��h;y�h^B�R↥-�m<��D�Ș|�jRV D��w�L>E����N܂H�!Uh��P��e?�+�f&�J�0Qt:���@�ˊ��r�Rb9-T�4�`�[?
��(mO�ɩTiƺ�m�5M�����q��ަ�h�&жF�Zd�1���AY#�j�J�ϳ� �����V��D��ૈ��)3r��""%�~�6��A����wλE�q�WIQ���']2������>1%%Aa������"�Y��(�/�Z���L�/�g�M@���l�(�x�́�K/�IX}1i��7��IyR{�i��"C�M��o�G)c0�B. ԭ�;>��Wȯv���yxNOP	7k󑑂��>w�i���@f����e����$�,���錁 �U:E7����c�SS�j���؇�ڙwo�<�=P*������n#�6֌������%��6��yP����QSK$� �i�$!���b1�w�׭����R�����m5��\h9ud�����k��+r�b��������GCm�'��/��KF�ఖ���
�
���iY����q  ��+�ÌF�n�
~�ּ9M���U]�^��-�f�<�3�C�"ؤ3]�QO?�h>C���4j�����dmS2s�uL�>���58-���A���x�����)Z(5�D�xO�l93�=�g�Y���$�޸Kp�驔&Լ=$��o�<��mzdɖ���Xǳt�[����0v�@�9����eYwO����f����y�1x�dev2�0��.���|���ϙo5���!�td�v�zR	D'�j�(�@S���f�5�O��5s~��7R��-;�-��03�5�3îΦ��g��©�Q5A�.m�r(��O�mr-q��R:ˈ
��N���	�� �i�C�$�,x,�n�N3Ax���˵��|���f�𡧋�d{�4X��w�a9Cs�^������G3��PQ�:��.j�M��xP�u��g��h�CJ'2}����6�v3��m[����;��-v�e��o��U� �W���Hd)���zz�ȾSc��J��p���&��P��|�'��E�Ӱ�D9��#Ӿ�Lp�դ�N������諎��zrFGm��H3R�������[�.��ݡ�uR'�3O���~�e��z�Gu>����6C��$}l�����a������dg�y�1�[`[�8�)(�(Pk��J�yʕ`q��H�8i�]�ǩ�s�[���-4�/�d��](�fa�oڥ��J���QbJ���D�_H���6�r0�|$�Ҍa������K�f�zrO=�$�I���)I�#e���S�I�IjQ>��	��B:�,I����Z�<�(���q�<�������� ڛa��住d0(ۃ�!.�����֔�W5�>q&�n���b��Ǡ�6�6�SY�(�����9��v��XN���ٹ� ��@>f3�a��P� 0�qj}]x�h���&��$�'h����k	�#K�|G�rmb�z(ڇ��R#�$$ )iO�;�	�:�p�:[�\�=��ߎ	�BR�-�n�I��`���dц�Or�as��3��>��JN��������8��=�'�˴V�T�̝�8H�?�����Ə�`|��N]��C��r���j��;��?�C���4� �j�'�q��Z\���ޠ3K䰇9Bg�?ٔ�!Ro�N#�ҋYӺ�%%ZmWM}��7gfx���F���EJw��,o��Z��4�ۈKt`팖��?�����jp��k�C`�#��I��{km�v�v�MN�5��bx+�Y��f�=j9��G��jG�l@\���c��h�첟��R;�,L������D�a�`���D�-�7�1j1k��e4S� ����0M�Ń)T�پ�/ۇ�R���Il�����TΘ�7���eq$�95�����J��H���b���F{+��0�k�9=�uiҺpD�����뫇'5����)�|Vԡ�Vc��ޡ��#�3�v�6���卵B��<�:����!���cz�G�טR3-�'T�d�:�al&�����1��bX��ɣ��RF�_��p��5j�w
`d2�gS�Vcŏ=��;��š�l/�����fMg�C˺���e��td��7�a�ZQ�J�-�^w��O��³�`.�7o�?�E���ٙy.��rG �T�4���q��hסɏk��[Kߒ�d$]t����-r!�*g!-_�jX4^Hw`H��c�x�&�#�A{�e2f��}��	�&���ƐЩDj��š\��`�=lP�p�6GO�bW6c!�3+t���cAB��MI6v]2v�'ȟ�����i�b�_��-|6q,��~i����~6]�鶞(��`/��J6<���?z����"Er��������;^d�� ��ƕ�B��nb��pocaq�p~�x�X����7ë��6�Sk#͍�I�JY�lޛn�� �BR�QM�����J�oE��:����6'����2���_�@����
p����=�6�"}ጐ*�r�K�:�MWUH[e��a��v�H.�CX�3Ύ��=0�nM�~��@��&�P(����͵	�Z�@��g�pX"	�|��	9�=����CH�aVB�uF9�-�v�y���觲�OndC���3��4���C�zV����݊h:\���'�	j	w�z��(b�{T}pgQ|��ӵ��C����h��7�z"2D(H5�'v��	��nĉ*����f�� ^��2��SW��in�P�&���"�z�S�����̃�ӖB�%y�5�=cI�1#{�ޜu�;f^̽��2M���p/��[?�DrX@��.kg�����v=[���`L?���L��5\���=����ǽ��,��uJ���;��=!�2��ژ&��@�ؓOV���)�60����hׯ����	Y����/�3�k��"�5{�?&�r�)ƨ���%avj*��2z�E��/ �ԉ3�bs�����v�q��(���z�t8u�`���G��Q,iP�H�,��<Npԫ�q������W��}( ��@�����X�̂FT�"��0�����~��4@t`��-O�Rj�f��[XG�R�3�};uZ*����Y��=�nWF/e�HRq��lA筏2y�1��6E4N���7�Xe���%�D���Za��[�Շz���Qn��5X]i��O��
��]`���������ĵ�/��<��t|�� �1勼��c*n]	q�)�٥�����u�8���B�U���w�R��VObvr�Mp_V���<�}����+gq,�~`�~{׮��aXqr˟���X�G-�@���L !���\]؄�������*B�no���(��'�׷�ϣ{�^|����%L����ȵD������:���Ҵ6���]"��	�����/�%��(��_A�h�/���9.����9�ǅ����R.̱�,Tk��cL�*�a(�6���uCD�	�D�Rd��1��o���x�܉�~� �m�X�%6�r�ɥ����lt�q^���Eh�ő�I:z�u��ԃc�1_����}�ǈ�Sr���;�e��!�%����g)9��"�gr$1�������ߥ��G��� ;j��y�S��B�**���ns5�
`�v�&�yN��@�	���S�!��~��J�qY�ȵq+�7�<Ez�|��t6��et-���}\�L�ܖ�	g�Eׅ�M���J�[fT�L�`�֢����6%4�G�l�Y��/`.������v%��M��)#��a�&c�]����`2Wr������kHO�AF��G�H�s����%���p���b)^�X1���kW -@�u��e��W�J�q{�B�4̋�����[�Zi�w�Z'V$0�/\���r�T�᷂[R�� �^i���:�n2��Fq��3X�ۮoR�� �I8�����i)=P,���K��ȵPs���g<��,�B'�~��RV>P���e��w�Nl�>FTK1b�B��:w�o�KY�݀qL<�o���s���<2m��H��,B�*��(ѫ��;k����R��Е�M���W�`����2妱�a�������=�k����ad�D���T�#�)L�Π�hO�*A2Ӟ�������+;�y�k�{~N�����o&� �*���pQ�EH
�ŭ���U��H��p���z��M�_�&�:��d��,��T [o���[�:,�h~C���v���g����k��A�@�냈~��;P�0/ð`*ş�vˀnԸ�\F)T��h�"�=�v������V`���Z��rZ,xF���q�VL���x��<+�o*?v�*���^�d����t�;4�x��1Ķrt9�%� ����Y��m�5`���s?m�+Bs|B���.Q�L�D�>��~�<��m�Bw�D��s�y�5e���@�D�/��g������m� (�	���d-�-�<s��fv{C�T�;٠�%Fp���F"]i���������2t��Sbp2L�&=��Tl<�]���ܧ�'������NU�q[����I�����&B������'Uh�� pְ5A��w����9c�s,�;� @��^���/֪2�%��$9�}�����������+Ϗ�dd�`������ِnb��~bJ��G��&�Ug�ɞQ45�kJ�&���-���j�]�{�DK�B:�y�����۫D#��z� gW{�nUh|��6�4� �ؿ��D~e�e�(_�����Ov�a�/�F�����R;i��C�uc~�^��<�%h����5�Q��N�E�i&�K��pr�>�mm�����ߨ���^{T=+{��(���,UMc�����h��������XO;$�qQ{�w�)�-�
w��PϽ��H��p�3V���q5��U��Lj2��t�*/��^H��ZS�^NZ��F~st�۽ѿYK8
P2\Օ��Z'V���g�o�o%��n�0r��q�[�K��л��.�=z���,�c&ZD����>�n3)ԃ��8'vt�Y@��W��0�-��_�v~�-(wJC�/o?������T��R|�B���Tm��\ui�ũ ;ۍ���'�	��x�#�����} G^-t	��]-�`_\��~v5lo�ЙGо�N�(<�`��P%���p�n��!�<��}ƿF�bfY�M���.�[	j��z�sm�I�����W*�"�/���ڙy� 33& %g�B9�/?��̅�Q`�{m�M3.%1x��K}m/��	��F]ĳ��@I�� ;�����8���/��aLb�������;:s�=9x����mr�����Q�!�y+׻!S�w�*�R����a�"���Zu$T���^ut
�3S�t���*Y��®��u��U�2�����2��坳Fj\�+������/�Q��x:Qjor�낗,�����tTV�^|�76:�]�$B~���ʙ����P�Q��1�����A,
�����&�����r4�d���w�����k�|>�M����VF���r�ns��#9�*'�k6*�)Z^-^GFڗD6��O1�|ױ:�T�xt���X�����N
?no��h�8�dZ�G���7e�m?�w`5M�pR3�N��d/�6��K|-��ߜ!(�b�@b�1�<u�t-�$��n��dC�y�(�79�w���#��<�tﱇ7B����R\�)PH���%&w��/"q�ht�wM6a��xv�T86�0���-c���:ǼJ�ZA,��Gc7��E6鼦~�iC�I�sc®��#c��p �9��� �NJi�c�Fae9f��Q�qōUO�?��C�O�U���<�P��GO���4�#0L��a��b�ot2v�d���Jã��.�*�RQ�4�tq�+��dq�0m*��Wqm���S� ��'��R�A
Y�y*�Z�ͷ�|�é�Qgo���:q 0?��p��>P�px�X�x�5���j��}~T���ҿ%�Ì`�V���_*��CRA(d�k0��`�Y�.<���|
	���#�^I�\(�b��!sL��s�����DAoѲ�V��ʭ��'y��q/���h"�|�Xu�ӌ�w���14��С��y�.a�������$kc8�"��wl��yL���N�i6m
�!�+�r�`��� ]J�����|&�4�?��(�l�a*xR��[lF	�0޷"�V��dv7,��K�iW��э��-��4	8�m�I�7�@�h&�M ���$nex+[��d��\�YD��cn|�|��ԡ��r���j��{��
Rr�(<5rnn$�7
����+�? �H��IK@�~�ǡ���Pe�.����R3��+��f�K����+�,f�b���E}Y�|G�h�߭�	�>�$y�}޵ɲ���Z�N�]��ʯF|���>UOb8�G�5����!�c�����8zR���*@��xjf>��#��/��+���x�S,��;Х�;�E��8!��q����P��N�L� �uϑ;3����*~.���EP��(�R��q=���'4��R���f�]���ݪzz�|C�3�c���+_�H��ݧ�3�9cl{~�8Tz���~�C�#���94�
1��w�*�J�KT��i״6� �u���l'�����*�ŏh0��{��k�)ViM�o��ޯ�6���wX`Y]�����X��R�"��i�KŲs��G�*���vl���q�ą��[YJ,�5EG�'�֮��HY�"7���N ��0��M�H%[qt�s<�qb~�%��H�����>G,�y;�ó�?'�n%3�+�����鈐��B�40N���=������5�8v��L�N��"#�$���a  ��
,�1�y�bD`��q�S<�(}俴N(]"��Zh�4��P��-|2�E��B���8�Y���z�S�-�5��)�Ƌq�x|��T�c�q1�ē��xP�[�߃�]�(�
��ܛ@�̅G�|�-�#�<_7����y+8�O}R�>2�2�?�.Ƈ�n�*��P���+W<�~)�9O���K�P�!�P{�G ����:�w��يp{�����Ü�a��n�J&F 幮�M�ɛYnF� yO1��nJ�
 �f�1:�qkZ$6\�KH�%�ܒhB����.���o������T'4�u�?FOf͝087őD�^H�~�^d����y�~I!!�i;�/�1�jp %��yN��
�u?��gx���fժt�2��ߨ�О�[�.I��3;u�+��r۵߱�/�')�����.���Cd�D	�gi��QG�]�1?�(� �%�3]Uy�0�
ǉyu���!��}Vۄ���[}��rs$Yw�q0�yl-x��+�ɨQ]���薂���M�<���� Lw[v�^#�w\&a�N����&�e,�j�;>�<.c�,;:*ϋ���
�q)=��.�X�[>$��Z/����rc���̜���ɼ�yj�~8���P��_�=��î�V��J\;ʠ/�_� �T����o��m�q�5���4Qd�5�c��_�����*�,}`���1E�ߔ���ә��������{	��A�9���B��l*�V|k�4��r�~�f��5������Ҕ��BLb���v�<Կ���t�^�0��:�=��/нѸ̷�*2v����x�c�e�ᗯ�#^M6UE����S�ٜ��j*b�I�a�2ɜ�3@��%�(^�2�5\z�����]�^K�4A.��v[Hj077AA:�\c+� �z�~����N��+����iHȩ�)�~wt�fL~�'��.c�Ly��mr�h��E��V�#i	��j��9���{:#��%�Q��kѡ$�S�5	�e��"ѡt�գ�lD�&�����S:�P`�W�),�ŋ�]�B�����C@>qK|�o�z
�N��`�d�kZ���Y<��~������H�KL/��	��~�KPt��۳�y��`���N����\[-�Q�K'<��R�����Ȁ�a����΅�6��-��rW�Q}�c�u粁SNӒ\X���kNS��h1�X�IP�I�4Rp�G�i�dl����H��߆I'�Xm;dp��*��B|ↁ-�.���٫L-p�9O�y��Q��A�#�ۊ�^���u1on�A�'�c����Q�MuG_e��+�+6~|m���p�q�H�p��]AL�b�R�*d����s���g��
���#\ \�Y�~��9�f�W�B��b�Q*{��b��YO�0!���\y�]K�+��ڝ� ��&r�F�X]�c��m~HpX���	��JC�I6�7ޤV.�u�gf���sZb�37XH��J��M�w^��c�TB�SΨ��m_CS�c�_9��y�������؟�-r������f����ă��қ lî_��D�u�[���s@�9�������N�������'X��a@k������MK�x6��>��4{�,=��W�d��E4qjR}#�V���j�OD�&�=��i�A�EI�����h�2��I��Lb�/����4G�	������\Pz��}��])h�ޡO�t��E��t)2��P<��ؽH`��"v���a���;���)]���{Ē.�Z��΂�����=����2�����h�;��6۱�
��
J��w,S
<���^K�����Vb�_�  �d��#/B�S3�`�,�6WI�)��ׂ��`�D����/D�ɭI���Y�/!��Y���Y�fa2A�q�{ɍ�^f;�Y�����L��d����3F�v����rWEk`d��X�u;�u	m���D5�O�TO���?��\�a�]�R;����C�Ut%�4Dwe+Ύ=@�
q��*`����~��G�+���eW�?�{�[d֒�9nA��֨�{fW]"��'HR�2Y鲙� ��̽���Fg�y�>���،.8��"��rZ�h�˅l;U\�}ݞ�ߘW��Vd��t��g���F�0e���tA%��ǰZ�ol���Y���!���`�'�u��m�>p�FE��0���%f�6�s �D�j,�H��PLT�R�C�`�@�m0�;�Q��/B�B�Xq�f
E�؎�Ğ�`A�	���$�����lZ��A��i0,�z�b����T��+�`"k�F򼸺���p�����TOi_(0�� �-�D΅mh$��X�-1��d8Am�����٤�������vlH��n2@BO'�O�5�W����Xt��vM s�8#�ю����k����<1Qj;|���v��9:D��FU"#�#B/#��rNM5XG�;�8%�i>N��ܛ�y��wUk
L��@^�Pv�׮���C!+h�x�%`Ŵ��_:���e+V�s��*�����Bˇ1V�⶟ta{)z��7Z1'������/"����28I�����Ƶ��漧�*�К]j���ݽ����U�B([U�&A׎�!VD<qxg�C؂=�%��M�3N�$�pƳs��A��7���ym1C��Wsn�)���83&�B�R�y;ő�>P#<K�K����\lD�4�@��Q`�&l4���K�j�d�y0�lagv��l���!	=F�k;�}wո_iT���=�X.z���=��	�5U� ���1��Æ�ݞBh��]��s1csz\�\L�_�9n�6�@?�E�K�sqhnV�C�<n�C.�<���� ^.P	�s�?�u�ط�X�E�f<�k.e!��%���7C�$�p���T]��!EW���H)��vIֻ7ݼ'Y��>�5�X�}�+�����z�i�e!�?��I%�Vg����v�@KZ�/x������;�^A��S1��g3����E�w9�VLo�U`��+���p]���4-�T)�-�����DQ���e�0w��u�ږ��f���5�c�~b�g*���x���3��f5<���f��4���/�" �|;C  s 3Vt�iEѱ�]��i�#鏵��f"�6ņ�����/9�RbL�=�;D	�a����CO4�������������F����{gQ.���� R���boY��
,!�z��̪7�BlK�����eͨ2x6�hg1�|���r�}/SA�8���(y��_6+m�]�>��9.rز�+_���Y�w7�+����G	�]��������4eN)�G��`=p��`�:OK����`����	q�S7��cy����n�\�@�_����`����	�����Z)����]����zd�"�����%�Pk���PЗ���	W^�gR}E>�fBm�=���_HB����C�j�D	�AŅDut��������H��sd�B�����)S5*l��,���l8S ��0��*��8
�lb:��! ���4�~RM��dl��=�ܩ{��̽�u)iD߂Z.&��g�7 ������<u�{12(Gq���4�5�&�6�K�
�����=̰���� �xu�����*L�2t�����m���G�V@+ú��ŋa��Qz>�`�����Ae/Lƚ�-pz{��d�)��y Ɛ_s���U��.~�*5.+�������ۨ�8�~d�ω�_�[�%%l�	{�aj3��5���J�0 �ǽ�"�i��NC>�zD�3PϞ��k��qQ��!D����p��!GOpP�G�*.\{�h�9c;K��Ԅ\��xo��0˥y*܅bUL���6ͼ;�ՠ�ʁ�\'C�d�=p6Â�읃���c	�_F%nnQ��y�o�G�tbB�Lvia��o�Z��J�"�ÚȻځ�qgׂt³�2O�&�:���@�NA@x6<R��sU׈MK)�%yM�C���5�Uў���R�m����z�5vdXxQu:���c�c��R�]���pd��#���I�_?�{��(9���WoR"�;��ƛ�"�v��U�)��ב:|e��V�<��y����B}完��E�7}��:��T3�yr)�J?-Q����&�`PH���`�	<���,�PŔ<�7*Z[	�(�^N�ڟ��~����m8#���S>���N�٣��3��� ���:ʱ���=�N�����5Ǫ'�ʩ���-��v�
�/%�{�;Y�Nc��v�K���"�.�7�sYsׁs�>�Gָx�]2�.T��� 7w�H��=5>�������w��g'��͏�A`�\��`�	/�����&��@z(�7���	��N���1�ٹ�Sڙ����%f�00 �Q�G۸-낹��=�h��\�E���0{��vs��V]�i%4������8�?v8���?{wT  *m�N�JS5灑����MW!����Kd�{Ճ�(��0.<u���F<���a6�� ����6���ɕT>t�q�!r�2�_��v#d]�uˌ��44���^mž�����b#�1�N��= �.ԗ/�P���:�e��{�]#1�i�\O�K_�=oش��mu޽8�u|/s�]Q0�*oC��A��r��VE-pxPd�(W�@�$���OT������I�u?2�5��C��&;���rQ�XD�s�F�l�c=c7E�W 0-]!����
����KU���`��ݷ�$�Rf���{Z�_|x@��پG�h�.ȗ}�t��8f[cĬ�uϠ(�I-P�3���mM%T�@�P��-_}Θ�`��=�X� 8*Ǖ�����4ے�O�����R;�O���kZ�E�M;Ǐ����k�z�Z��7�Q'�8*5��'_�y>����n��h�4�ǆ��@R`�q63�´�����<�}M
�Ț�ڳ�U{�!}��h,%u�}@�u�ԠBʶ��y�֘,�H�]�9�=�
�բ��0
QQ�!�GIL֜�ޡh'�c�U���@���E�<��,z��}d���J�&���qY��
W�qT�[Į���H3XZ8Xp�U�i�����b���g=Dт���H����j9Q:tx>d���p����u,��.ܴ�Q�����H���yE��J�(*�������R�J�^O^4zu�¨�^�t,N�+�=�� �S�j`|�:�{?~�GV�'��-�w��Ҽ.wU�hϰ�R���w�+y�H���ҫ��B1��+╫K���,s�e)�ᔖ~���V��+��L'��E&ݦgpt�<���,[��(,Y�Z��/�F$�V��:[2��Y7��3O�(������W9 ���+
0bm��
�(.=l߉�3j�zW@��z����*�z�.����'ޭ��B7LG`�=H�O*Z �:�7�qNoZ�V\���@�3�M;u�6
�SǏ�)��3	ޭ���n��Qfe	�䔸{Y3�@�$��g4���nIՎ>}b����ۺ{�� �DƑ��������^H�x�\'��C8نz�d.l^H5���j�Xv(����_Bo�ش����&2N�� �.�4�o,���C����]�oOD!4��2��r%;}�y/1'tS�]0�ts��a�� LC[�)�Y"-���3v�G<�_}�*�U��c2��CL����r��-�J�r��?�ۚ2�Ze��I`e[�����}� Sf�q�kO���]� ����1o=����|Xd+/���kbr�H݌�����z3���,A����by�{f/�v̖x3����
aIL���FZ����0=�3��T�H9����S $����-��K�m���ѫS�ՠ��)���%����#��ߞ��v�k��&���Fr�'��3Q��%U4�״99��9º7�tMW����y�\�(�\�%i��M"K�"9�'�秪�f	7�'���dM��<�⡬���sS/~��
 Ǌ�ޑ"E�dAr��O��s�$z���M+���I��EG��0^<�UCު�i(�j`z\� �O�n�<nw�}KS��u4B��RWm!�:I��x�����i�ޝ��a���.��9�?�T ��5�gR�/xd��F��U(�݉�)
�Zb���F���N0P��/��>����2����ta���hVǦqPU���NP�d�x��2,P����:��b`��G�4�I�>��1/��8�z$śE=)%��,��`�Zg�m�|efh��T{�a�1*���M��?d,��Ǥ��6��b��DZZ�ad��O{��Y���|C�'ΐ�6��8��F��s��%��By�����{��6<`���0q�� tI	1�p4�i*v`;߭�K��?��CO��H �K+�8_���hG�V��*�MNz!���-#��d���'h��!\]�1,1��1��3�"l�f�W2�,� �ƽ��] ���^�(���
��M� �c�˝�->�M�~Q���gު[_Q�ɢ�L���IO�`��K�����]�v� �ꖨ������b]꾯�/��W������!Af���������ny^�,��dK����b��ֹH���@*<a*�X�]���䇚��������yx�i؆l�����| �
�PY@�{f���1����'.
3q[�z��^�m*���s�Y������}��/lI�g$�	��!���� Sr�=��5!V?Y�?��yhq���f�=#�5@v�=A�~}S�)��%�`��QŌ�_g��|gH �� �i��1�Lc[��a��k���z���0 �� |���3*�����]T�a��g���uN�QV�0\*�u�ɷ���&�y��=%���Wr9kn�**vQ+;��r	q�����5P/c �}	���Dq�:>��Dbe<�Z�%�X�p���IV��a���5�Զ;&��ݸ �F�>S�q��{oZau�V��@����;\�B�
���>QgZ�<23:�	��7f�����V����$�Ku�+Y�I�m�ӣ20���4����!*?�٭<5��*�d�b���4O�?�-Ϸ8_��T�+�����!g���a����8����`�y��'�,��hD�lg瓄�8�r�o���^C̀z�� 5�=�ků� ��u��24Σ�m�9��h'u��4�B�Bo9�SL~!FW�+��Հ�;0��?Ȳ��H�s��s½m� 
>�����
Ɣź���\GߟZ�ΒcB-p4	���ߋgG��pH%#�/�K18�o͋��� �����j��7�< �ׂ���PO���WK�A�d�"=/P����[�R�܄z�k�U}7�̛��gI��6R�%$#�b˃��x��Y�P��,�]�gKj0ͭ[����cY8b�,���H?�r�s��M�u]"�5����L=G��|%��렿S�hZ80�_��h���o��Uz��^��c�4�y�U�����*��TDg�~Ԋ��8P�F7�Q!�$�{�M�M��!���]6����es.,|m��L ��(2n׶�e�X���U�M|�� ��5䁂d�u��p-�Ȭؑ����J��M�6c��#��̓����X��п��8א�6º���@F;E�\���� �hj1���?�& P��
��O�bT�]}�wvS�����m��t_'��!o���$֠y`;���	�͜}�^in��fw���{�h���Cm���PII� c6������v_5�xZ�C"�B�O�=G����u�2H���ĸ�ۓ�P���EcE+a��L������P�W�y��!;�s�~�<QdH��x>�M�?����>�%i���W��r�u� �F�e�]���?8��:o4���E^����`�O��X�(�Ct���G��
���'�����Փ��Y�r�xCB6J>x.�ҕ
Y!��4>��}aU��,�5h�ϱ�6.������.����ќUŊ�I��S�/������nQk��)0~pΧoa�pc�?�b�Ϲ�pO�wy������BC��j��S�BK�l2�t�(��Wv��jW���^��ݚ�ؑ����F#�,���0*�6�FT�t�!�\�R{�I����M�꧄�[��'>ɻ�vG���Ǿ�x�5^�<��̓�3��u�b�
��*	܌��R�ʶ��~<��.i������dI������z�<�� �,� �5K��沬��2ؘP�	��ټ�'|��{R��{ ';wl`�r�=�Y'�"��K��,^�������`y�[]u�od �PktͶŝ������=p��S����yt�we
���:C8�dg�K�19�/��@ƪ��=..�h�T6l!е��Q!��a�����j���|�ʆ�]7��4M�tbe�M��Bn� �<xbЪ�Nӣf��N��F:$6p!�Lp����ٓU�:׈�rD3�Z�r�C8������+UE�fY�i��AJ�1�x�D��x9�@�ýGx���_XY	��A�R��R+1��e��)��= ����˰p v��Ё��V�g�t�������`���,��xF�<��Sy�|���䫣�byl��ďVld����P����G���j�}/��ڝ����G7�k�F0kK��kSn��;:�^���9#��:����w8wk5pϤ0tc�"2`l�/���t'�(��ߌ�Vu�tgn��fi )󢅒��e�[���[�K���`�{q=��W ���?����%,A�S�l��EO6*�Hy#��6QS�(�H8�[t3���bPԤo�~����j4�U��θ�����a�ZP/ei�eww5u�}�g`�b�ș��'���DM�?��G7q�%����jV�Ţ	�!_66�F��j�Y#��;���O������lY�Q��?-aGx�w�T�4�/��~8�N�u��א!ߵ�![KG!�6?d��#�<��%�=^ËQ�`�쁱Վ˂�)�(�7��]C�)m#�E���U+N\�s���) �G�OWrm��}:U���}���نZboV/I���c9M�xI�#�����ߚ�d��7�W�&�_^C*���cRLȥ��j��+ܰ��(��'��ae��mU�J�a�=���X,�����.0ڈ��5��6�5p�Ϩ�N
��"SY�BV�s��X�*~�"z$�x�_F�FU6H�:���{q��$QU���e�Z
s�h�$9I4*�到6(�f�>�8Y� ɞ#��֨)��҄�f@+�>�?���g��U��rzji"0������^ɠ��QgUR���B&^x������V3b��c˞�=���NR�ӻ��<��Y �*�%��������q��9����kF��K-%�H�qy��$���(^w����"��#~���[Ԋ׃�3	H�W�`s�n��2�t�G�:N{>fI���:V?�;�Y�E꨽��aN�W7�T�FZ�p2�� y\-y�1�@bc�e\e{�Sn6�i��S\�)�r��ǌen�
�I%<^9P���.��5e�Uqa/Až"��4��]��/�o#�Ｍ1�(A^Z��?u��P�{/��Q:�p��Bn�X��R7,��x��d\������.��zj���>�>��[e0�%��};vy�z�3���n�L����+{U�ڸs���Y��־@��|d���dk�v�:̧��k�vg9ק䀬uY/A���)P"�@��DY�`�{[��Nv��s{Z���в�1zYĄ��q�ɑHl�	�vH�ɫ�j>F|=���`��JB�MsU����Վsz,Ť5.����mz�����5�p���a�n&K��,͑��̖��B�ןhD�MXE+�8$�Y�A��AwT���	�X�i�($�/L��4w,߀� �˙b�E����Ր�5��468{���e��DO��U�G�+��(��'�6��ԏ/4;����ۘ��Ei�! ��qd����)j��{�KbP��X��4�$�˯9����� Ba6暣�����'A|��4� 舧�o7T��C�)��Ln���o_Ej��F����� +�߭����J��Qd6l�Y�]G6������U� ���L�D�ly���+���	��]���KfQ�����.*�h\�w>��>�Y�M�v҃�A�w�%���c�՟�*C.��mm4�um����F�Wk;'kNғ�-�G���ch�գ �^C׉V����v[ʔ���1+���X�ct��a	�ƹ�[lH���n�u��|�x�F�*�!����{'�@��ĵ���ϼ)v<q���vSY�"m2G�G�㒝"ls�N���G�=�@c�fe[D���l���
^&�X�1k�7~I�ijmE���*ʙE����
D���¾��N�h�盤�)ኛ��򚞎)�T��=tu��I���#lhn)Ӝ�k�gP;��M(ǡ;u����pMF��u�FJ��gXBK拐��0���2KZ���	iBO�xX ���w��"��=�[B2jo��t���?�N:��Inb�L���*��|�F�C�*no���:�@@�2���3J	���叔��A�}+o�|���?m��^C_hS4B��z/+ϠIC��Z�ݍ�ژPͺ��V�Q
�1��^�>�o%�J�\�_��k��]�k�f�O��+?ss�?��&�h �-�w[�Y�YN�DE;��qO�ib�����xc��c���D�wd�v��voc{1Q��d� y"޼��F�������>��UX��#d���*�d���n�Mf+��{���,Կ�0~+��qͫ5�)ţ~O��)v���T�LU0R���Đ8��b�YB\��u:Ql�#D�i%*��(�WG���(����:�lc_�#� ���K63��/���������������̃XHٝU1�@x�]�'�.uٓ�E*`�ʡ	-2�t�N�߈�wlP�/��t�Bc	�a/|zB�1w���ؙr�%��=�	PO؄�s�S��%����3g��}�t\�#0�)~k�s��oU����R���� �� J�f,���FQ���U��5�'�܉ }�(ONmH��}ԇ��#w^�t�e�Z�T��	_��[l�Y
�L�k�j▩~��#�|�B�}p�4���c�z2�����|��EQʈ�t�Uy�t�T��8��_+��Jqn��,]�T���{pf�:�_'�jӉeB�^�YÇ��{L�OIN�l�厢D�o�rN��K�%F�נ�m�:������KW/n�|��	o��]����,Pks8�0��Ăd.u�R%���W�H��9����G��H�(\ðq."_(+��*g}" �R";��9�\�]ru���\FA��~����j�lVݹ&6�
#�_�X0<����@;�������Y�2�|���������;̼�1�J�a�<M R�0�Z�O�be�k1�똏�%�@���[K�J�������!̼̬�g��v[��%}�]��Q���*o����%9^�D�����C�&l�9(�#s�31��tp.7s�ڪ�wي�Y\��{����=)�J	�o��6B��	��@*1�1?�!2^͑s������7H��x�xkw��h����R�{��B�K����>p`D!�@�Z�	�u�q%��ш�����N���U��ŀ��*C|.c��r��<n�.�<����ڨ���z�K���.��Yc�����|�M*�u,C]ڶF�
�Ua��Pc���/V
E{���$�r�6�#��נTr�BK�~a�Ѩ\��31�q���L>�� �a��\4t3Y��1��x�M��Y,�l֩�8�u؞�-�Ho�!x�mx�	V{*��>-�'�"J��n���n1����Z���훸~�bA�B�^��mCG����`U�=*0s���f���db�c�$�$h}�s�ړۋ�T����υQ���h�Sx-=���~'�?�����t�Rǫ�fEB]�.�,����@���e���fsQuj/��-޼a����ۯ��J��]�n+zcIv!|m�sZ�9=�Cw�g,O�����9a�.e�xP�f������!A+���S��b����z-�}��r���0IN��eH 4߅�&at�	檪s�9�KЫCV�����8n�&������{������5��1��䶼([�W��f�M{j�
{K���x�ws�.����	Y�m�-�0�b����ݒIE���u⽕�`;#���W���J�a��⑟T�y���H'��A�CQP.#�៸�Ɛ;GF?Fƥ��!�dn-�V��N�� �L|��]��g�3�&=j���G2��<n��R��FdU x����z.}R������4��}��B���k3�����1�g�[��:���m����u���
ɢ�z�U�×�G��R�Tp��5��w��Y9E��7L�����ζE�yB"��WIȾ<��	���$@�|c�ֽ7~_;d̀���b��׭�@���<��CW��]�<H~�����Ʒ]���:����+�V�mΛ��m~��;㐘������9���A�����j�uR V�oU�	�ɨrw��R�O(�����0nQT������*cL��\���T �<>s-)����a ��S?xK8Q�&��M=�_�����]_h|>G����M�0Q�F�GѳO���\�*}:��pb����6Z~��ޤ�J'1�#	<`����{%�ʜl�Y_K�Ⴚ����-��� o������dҲWi�컕j.0������	��Si�2�!��� j�i3�r?]"mv�mb��)�;%^u�Q[vRb�)Qx
쐋~>�18>zf�3��G00j�d��i��%U{��`���{��%����qq&���Wjn�����O��̵�����<o!T����C%�h�%W[V�Q����R"��'��`Z�¼���P���x��{�������j�Ɖ����^Я���z%[��ӱE*j��FfSh��R�Ǆ�r��>Iy�m�"�=�[W�*%�\�L��$���D,�¬��Ҍ�$@��K���u$�������	���
n=
���C����Z��_&84����c�X�����>.�*d�Y�G�Y� Q=��n)<ݠH��V�U��O���G�bNѬ�
ťN�CI,�@6�9�]�S�+CɌB�8,���[�.Kl^�Ћ�#�J�w	��݂�X��_�vր���w9�5㵃��a����=��$�u����x~n�A��>F5ԡ�~Ə�B���5��<=��-b�GkTO{�n3� ���.r6��'�TP֓�".Ã�`���^����X9�U�d6�OK��:�Q5�Q�_����e�HpF�]�}���J��<��ꏩ7%���͢RM�ze :�c5���m�/b~_M���U�l�8S����98Z���O���_�����&�gEƦЁ�-� ����7y$�a����<�?Td�#d`��QB~Rk�h�"���ڌߌV�^�9����>n.�B��9qI��^S��lk��������׏,E?\캲����,��_AŹ$��AvMT�V�(,�9��?Lhn Je������"_�$�K�ۿn�{s��4c~���Q��z�v�9������fz�|#|�`�!��hw/�M��2��G�]�Z�z����<�V�N�D̷ٯ�-�]�X�Q�Vד��,m��Z��#�bj��y�~�H�3i?�Eh�՗XW��A��w3�7��Ț .x%�M����ZC���>ij�]�U+�S��81M;�8E�����X�O��`��oA�{$����h �)J�+�	��
C���� �7��)�1 ǨN�:j`�J�|����NJЇ�.?9�L���lxR�>Rb��aN���>Ģ��Řix�����ؖR�!*V�_HR�v��_Y3J�K�S��������.������<z��W$�*ʗGL���d�O�
�xw��U_*�V�߼!�P�1��P�h��47I̺�G��M�o'�zm���w����U�F[�r��`����lx,��w�3��_8�0%��"���g�a�_���y&�6��*aQ�O;��C�׿p��B��;���S,�lw��ݳy&�{�ќ�s\, y�k��6{maL����'�e�ƈ~�X߬+����@� H����(����^S��-HvE�� '�Mk���u�߹�
�F���9;����
�Q�2�:��9^g�x�A9prM?�_�^Y�L?�%j�V���
�=������S*���=��6���Ra�����B.��n9Ǩ��y�m��L�꿮�����枤]�_��X����/�q"=��slBiT��^^�>���� 3b.�[�������M���� u7H[Ԅ0����D"B�P�I�����F�zH������ܟ!�H���$Q��S�yw%�4$�c�\t&�J����9?fc+��&cY@��#KۅS=�NԩaC��by���z���~*W���G��;Z�@y�5��ޡ'��q� �Nd��h�_BX*~}m��E�PI��p�^�/�+j�Z�Ez�a�g�
��yM�[D1�����;�g|�@���K�Vi�8� f�lA^d��ү�D�&�#Ŧ��۱|;�']v�7C~7�j�R5ng�_%�^��K��E�zC n��SI�3p���oEH@[���L��Wt�d|G�at�] �-��C��9��	/^bt��ĵE��m;l�ϙ�� n�85�X�Y���� �}�#�a�-��MM�)d5&W���fV�b���rbPR���qc���2���Ol�a
�L�_�e�R�ʓ�h_м�=���j���j4M��eDg�d�eGgM�TzH�k}��3������}��b7t-s��9k��f�ѵ�����E��t�-o�}97/����Da����7�����U�Bx�7�����3Մ��ԩV�Xb��V���pU&����� j�ۘ���N����N���n2X�QD�{����Y�8<뼦�%� ��d	�9lZj(������2���m�i�Ag����,� z��I�!^�1'��9�r�*��L��G+-�e��u�|Hwũ������{6M��]zH���d�t�r�ψ��nm5��9<��L݄ƚg�%.[6]ḭ|�@�4��@=�l�h؋�
�;o�� .9O��I��Z��N�D�G+�)�Fq\Mܦe�(�"��Mi{O1�pǤ��m��BP�;�5�B�	�E�#0P-D���T�"�$���4�
��_Bx&���H�ǜ�%=�&��0V��.�Q"���xG,� C2Έ��RqA�.W=����łr������ 
��f�v���(���N�Q�C`����at��{����P|�:m�o�/�������킩��f��f����I���JR��a�����s�>��r�ɺC� �ҩ���['f$�Z�ALw|c"�9Q��4�5��wS��S���L�h��3���{���@O��Ϊ�b����|�A��%���4�'��w��/[^X�����xj����6J��`��yf�笗�G���rf�{��e�>�H�N.�9�_��+�?����Z�����=ps�����Q75�x�meF�4-��%�.���H��/��MX�/d��Ģ�:�8|]���;׺U��"|����S8M$
��I�����)��I�fa�>(�l��R���Λ{���#��z]��uf^��K���v���jP�Q ���`Cŋ�O�%1@:^^Y��2zW�9�4U��"�t9i�ǲ�@�R�����J���΃�Γ��O�.j�9�W�z���6�m-ʓ�s��m���Vo�
�N���g*�6A�	��m�Rڊ���,�_.�܎�n�1��o�! ����C�7�wR-C��W�~�)א�S1L��g���?���[�v�(�p�������9��n�BKܠ�1��,?�+)qk&�ۤ�V�[����ڍ�&��T��[�p��Yj={~����%�x�<��M�����������<�{����96�X�h���X} W��A�����ㅦ�����9/Y�A��eE�6��S����!�j
5��o���ҟ���?��l��5�CŶ�y8�$?PsёD�L��"���b��*&n��ӆ���ce4���6���������m��"���V�p������X���wmSbY����{ݷ��7�~�в�
�nJccU;�F��ß44��l���w�&>�Yl0�;��Ph��O(���uj��~zv�g�4I��FKEq]��zh2�<�!��K���H��\VE�pG����]��5k�������dY�"�B���,ۃ13Ĭ�g���# �]�A�ܱ"�x����b�m	)��ew�?��h#�8��n'?�9vu�e��.i�R'E��� t�~��M+g5E�/}�	-%����Оw ��=�?��H'`V��$Vte����4�1�M��Vo�:�y�uP��4��/�o�}�ʷ�
�.���o�>�{��h���8*Ἇ�C.�o��}�T��nϧ/Pԩ�>��ֆ"U=�E:ls�LEÆX��<6W��K�T�]7�n�\ܔ�A�DG^�ʟq�;�[/�IlJ2H1�vSg��)h�i���o��9����x,���,i�u��:[]"y*J��O�*�$�H.�^B���bMl���|D�O4~�96���o��fsXr����sMe���
�30֔��G�)���'�2J>Ѥ���ଡ଼���C�:n��T �1�<M����鬶�L�!z�l#e�e	S�ן(6�jՎ�}q)J��Xk�a��x�����m���<#��k�ϻ���^.��DA��?i}���Mr�(�[�f�o.�=W���0�՝�U�I�@�O��_;g�pV���+O\\Z�W�\�)d����~����a� cfe�%�|T+���c�\Z�<�,lb3i+r����B�mVkb��CY���Vb垨5˫0:����b�*4i��;�D[G��p�5��n)�?��������H'rQ	���af�b�㆝��_�t-d]��;�/���[;�,�u�6{���Qp��C�����˿!��	(���)��`�}A{`�O�F=dX�O��/3$!���3<�]W���sv#!�j�
x����v~�pv����D5T�Y1��<���>�L)�pGiJ�!r�U3��(��T���}SU����4�Z��uӉd�%O2%95]�z��;@4D�or~��/�jg�ʺ�%,�H�*��I��X�G�ѽs ���r9*�P��7�S`O���Ã�~w�N���\�cz����-Ylf;@�=����ip���ʛ'��Ĥ�!���<D�u�K؅�{�n?�Y��Xts��Ky�6��O��^�&K��u���hW�e?X;/u``Y�ט��D�h>�P+�N'�!�0�φ*��&�׃ ��a`HeYK��1�3!M袰����(�I6��&Ǩ({�.�� ��1&�~�F!҄���`��uζH�LD�T�~+=jv_&�-!�O�w2���%�FD�D3�����|,��2P��	\�}<�d��|���,�K�oW<���K':QϘ\,�Y�r���j���������\^�>�)�6�$YZ}�v����n��wK����1z��^�l����*����ej+LM�c����;�7�̾������% ����^�Z�oZ�C	*��(�|���p%0���O��lji�k�@�:BYݥ3h�NCuk����O���b΂׊5*�I_X]���
>�uj��C{�T���"���-���'Ҙ���	���&�MHz��[��4W���?�i!��۪G0��s ���aOf�L����&*
	�������CJC�B�B��j	Z�
߼��Q�r�_�dϹ�b���F��� ��t�˱�s��,}���U"Y����K��G��lu���,1� 9����KF�)f�o��}�׳��ͦ�v����}}'|O�JE��px����2?��_=i󇤃N9�w�'�N��c/��{�bP3Fߨ�d�����f���+��Q�}Pƃ�4�r��q{�`�F��a���5�����+B�����ڞ������%q�.@��9L�x�t�� ��I��5~X��g�b�7H�>9��F�ck����AMo�s�c���ި���Z���p������^�ӳ]7���� h��6�l�?�+9V9�^�)�)�1�Z��e"�-)\{~��&m��?a���;��`�֟j����)a����檮��YO�2�ރ�L�]9x1tn18@�(	v>��֚��X��U䴙a�������T�/9��`�+������GOQ��ӟI��Ւ�g.ė����G*l�@�^r�EԈt��`bN;�լC�����_���n#�Pv��8��ֶ���Qn�E���S3n�(n�w��Ȕ��l���2�����0f�F�S�ˤ�"E#@,�	��̃A��%ۆ|eg皽q�v�h$>���{T��=߬�=�*���,}�u4��^����rC��ש;�ԎM�wІ�x���ź����.]�����F�Ԧ��W���A&p��uB���W��f��"�n�ɕK]	�*R00���p�{��Q�~B:��/�ċ�q*�U�����s��FQK]�<WW���>���Fg�3D�:I����3��;U�0�^�=-'.@"�F��WE�dT�\�V).��I�8q&�(����-I��<��߂���[Y�r�6+����Ҟ��q���F��b�i�73(�c��{�u,�6_y�A���*�ڋ+������J��8>�ѷ�>x�B�(�A��_��8���]K�z��-�&��c$��K��1�8`�"Y��8aG�Si�K�A?<���)En��|������U�'e�Xp�VV��׳|̯f=���*�D�F0�7k���C���oZg�1	�C,���g@�P�ǧ���b���eQ͜��=�-�����偞���%�(#�p�I��}�6��.���!��X�z)(Kkʯcq�[4u��0-Ye�l�:�4��� �	��>�\!��l��α����=Z�{�K�63���,I�N���)��TBr����羧��G5�
]d"|��)kj��k�&����]����L�O+״��= ���T\�l��)=���s�ד	;As�c"q���qY�L&W���ڨǢ��ۓ����NAB��:l�ݙ���B>2�����P!��#QW�VON_��|��8�O[�;�;*U�,����3Z�uC����Gd5��	�%���V��Ý�0~.�0W4';�~y����6�mKų8��)��	uHJ؁��-{bX�17`%�?�F�I]�C�w��_5���2fI�BG�� ���X�%[�e�B��Έr��6RW�^q9���6o�v��U%�.צ���K�D4�}l;o�X���6�9EN��]
v��W6��EIB�#6|Pw�uJϹ���O��6AWk�V�%��w���T�6�CQ��PTs�+�dX�xZ:L�=Q'����qI^ mj�?r.�����K|c��3<6���Hb��/��*[�W G�x4������ݎQ�Tξ�܈�Ffٟq���z�(XV�-�����,��A\n����3��&#�(�4��P|�p�:�mc�x�q�][�=d�2X�C퓺�D
�����^�y�LlR�:$mYQH����E���4k����� G9܉m�FZKD+�6▤ �0	�J���g&�)oGT5��+5D�J\&�1�="�����KN�r޽m5�RRI3����1R�������F��YBx��]�%�_&����ń+%���0r�:�6�@C7�f�������R�ԋY]{a9����z��b�!Б�^w��{a���0	J�O��)�R� (_�[�N�&͚q����kۘxYdr %�o�#L�AK�3����e X��¥)�F�q:S�#�)��a4�Nr�����ʃՙ�7��#^i�C����P��K�V�l��m�j=�(�x�[&ܞ:cy��6��&h%#�Ԋ*e���� �1<^���!o�E�n���üW �x��2�=��X_R�p
:�Q��7Q�kH9�?��/�z���
A Mt�����O�2
�XP*s��t2~�U�9%|�m� �mh��xb�ꑕ9t�Ms�w��kI��"��=�t�dK�l�;=��������U����g���koɳ{K��I�O~ew�^�����ur?��As��-|#�����x<��~i��d���y�[���P�1�ܭ������^�:��W��+�^vnM�Q�)�����}�p��4c�<�-���q�HxP�t�����}�W�x���$
�'58aw�;�NO�:{�:E����zFo&:+�9�.F����L-h�_xz��p�R`����=��PU!�:�at]�.#���#?	� �R�v���5�� ���2��!�@�@lǇ�[v6���㤟���J�@����:eS��&���0י�b{��OA��`r�iK0,�5K�DA�ћumD�44��Dg��rCY$�����=���kQ����� )����D�:GW>���#Z�jaXȇ�k�wn�w}qm��B.��m����.����4�zv`(��V=�}�7u_s\zf��r0� d��>�!.�*�!]M7I��}����!H�,L2Ǿ|
]�V��]�N����*y��F��v"9�O��Jj��"|=�źO'RH����|����7kn;d�U58ӊF�]Q�m�P98g� l���)�<����r��<�L�h��E<XS�w�i�=�.:�(��)���In�|Mr'�u�"��[ܼ;�ۉ�dAD��5أG!
49�|����ɺ��M���f�z�[�`���zr�M���v����d�CRX�	-L1M�Tr0�	��g̜¼�q8��b:-�}K�X䫡e���Nq�����ᐾ��/�Hi��wh|�����E��6(�e�G2��M�=�i��^�!�,�Iۛ<��`�;[�'9�����֙����뀋���چ&s�%|K$��&�w	%(ʇ5�����!_9߇����q¤��e ���vcj�h���`�@1=�7�"�R�nb;���%�|�k�Iڭ�zyߛ�𸛀ˬ�;*��D�$'�:^z��E)8l�N��@=����p�7t�V����	1DB`�/��d�vlGm	�� ���7�K�~������l�	A�i��f��/~^=%H�0�ia�q���	�z���)�q| ����#����6�Q_Q���h٥6�z�)���c�1��u�zɺ<J��O9���e�9Z�?ڼ�df���['�	����^���4'����w�y��~�� �
U&��!q2�H�+��:3u�ag���� ��0��u}w�R�е��pp�D�&���{�����X�I���=;����)ƥ�{?��v�K�L|b�o(s���\� śb��Y ,^eQ¢�2�i.\ʦ�[ON�r	���s_�\��Z���Nʶ�j���Ҫr�b�4�po�)�_�������l�FdAJ���N٢
i��=L��nt���9Yd,c�x�E�ܽ��c�e�[Ä�BOKNJ��iZ\���ST����B��_Q�m�$UfI��^7�fx��
`��|�X���F�[ҟ%�o�8$1)Daө]�J��7�0���U	ڒ ��wl��������1�k��L�}��7N�R�]���Vq�)���B+T!'��0�p�ZD��\{[��V���G+ox��y|�����ۤ4�|��|�_��݁��Tq䞭�Z����u��� �-���0��L�n�Z`���r��a|04H֛*�=��=�k��{����$'t���(w����^;�GO�I�n&�Ms��!r7z�#�$� ٩8��������ߝ9��e�s�mS��#7���Sg����"S>K��aR�D0#���R%�>"������1N�B^����S��M,b� �0k޴�N�
���9����wd}��m�/
�sze���G�JF]}=5�Y+;��w��g�Y{�x/�;0��	!|�*�u�G8��2Y�0��U6��{w�w���;�%~���@%0��'=8�[X>�3z��<�m0��J	���X),Y��w��ie�����s�H�z`ۛV�E�j.�f���2H�Ռ���?O����a�,�S5
�C ��������A��l���f�$,��6�ɥ��jN�}����@�,K��7`K]�C����'Lbs8������D�C����?)��Q"�X�ҳ
ߞW��������
��o~LIe�B1Z!v]'L�p^��b�#��@me���\ͯ���$?����%D^��[��@aQ�+��Q���{�y@�WOr�|V�85� ۙ,=e��p� �Vk�d6�����J�®��uZf��s=bZ�X	fT.LO�����>-��	��Qf�6�+2`�i@����T0a�x�]1�K�����jem�
&�m�fHWݠA�Li'��Zx��O/�f���,�`�K�\��������>m�{�-��F訉 ⱇ6��>PK��wb�K<y�r~����i��c���^Σ��
�'�(�iQ��:������?r/�A���{u�st��W|ɣ�[C�;��>s�]:�e�X����I�I�3a�Wi����{p��ꉏ�����S~�0�3現NJ�9�8�|g1�ϫ�n��(�M��Ԡ�57~L��L.~N�9H���Z�a`��G�=���ލ~\���D�60��M{Z�/�&�bZ�i{E�hȐ>)f)n6z��$��J��%����e�����-'"�'�����Ϧ�Δ�O{jUи֜�Y�r6"ͩ;�U�c.��}�I�Q_bǊ6d}�Y�*6������[���?Mٹ(�վ� C(�6vI�� F���i�G��n!��Bm�=Cu2*���*&�_|�:��ۻ�r�<�/GH68��2M�M�j��8![@`��l]�-3�����ꓸ��>ɀ}t5�p���	]����|ͩw���Ⅳ|z�ͯ��\"a����D��$����29���{�7VK��q\�|P`����9T[J��*T���M�٭���da�L���8q������
L�Dϧ�ѩ���܎l~�m�~���J��#��z�����E��D#�}@4�'6o<�a�=h��o��ӓmg��+)�d��ERb�Ř��H�vş���@)#��D��f���e�{�&�����H[T:�S��Q��&���U��O��wL.>I�؍��'np��Z�N�P��s��jj������θ^z�A�oD!j�Q-�S���
]Bnu���F���+D,��>���3�j��[��ֹ8@����7�7�p��?���]�FBM5�*������easHZʦ|���n��m���٤�+�b���Sݼ�!��B%�oD�����TBMTQ�edt���/d��?f �m83��a����Ov�d;���u��l�����,��"������;���Lt�1*�H݀�g�v���HO�[ue} �1I�8�Ip�h��zBȕ��B&�C�v���/-F��TGg�)X�具��4��>�"З���x~G.��ˉ�P�dXHQn�_R��1�i�r3⼶�D�jP|��z�1�j����ք����Hp)��i�F�][�6w�mߘ��Q��l�6��gG}��f1��s��O����3��2�7E�3�1���-�駥��$�Tzpȧ��:P#5�)�h�hM+̔�|�L ��LB@��d��:p E���P͏Cq7Ȍ�1à����A�T��F�����#0x��5�Ӄn��gG��IUӸ�BΙg���/.����{�΢�̷J�,�"���{�5����@3�������Ռ�S`�P}[v�f���.�ΞM���*��5��0"(�?�]ԗ�hnߨ�_,�0�W-&WS�5c��j������U�p�$�u��Ϯȫ�BQ�}vJ힗T�#x�.��h6pg�����%�?*�C_��.���N��/WTD<ے}@��
O��>t���|�f��̴�~rx2�����D����K��]?3:>C~M���>ofGT��~�Ɖj�S{BQ�M}�a;�����,.	���t��g�S.�QZ^�Gsp14$��ɔ�}>�$#����.v>4�&����
�<
D���� �v��6�f�n�\��C��ݵ���׌ִ�@>�������M�-�afTP1��dH._�N��80)���!8�EL�����veAIC��J3�!����s�#g�9cg3K8�A�!u�M�pA�{��4��p�u\�n�Ob	r�����ǰ���M��:�>�`gqY��΁�鶂S��UNH�B�@G�)�:x�bE3�ڀ�M���$�JՎ�з-��X]����>�	֖���e�%o�5����E�r����9��`$4���Ohxc]HI���N|�>2��h˙Ć�N�k@�/
�#��uP�'�g��\1���)<���A����O�8��Hi.:Ň\E��`	`�U�O2��x�d7���gD��|�狵�b���LVؑ�k7x8��,��?\n�Y� #G>A��E�^̓Z���d�bG"P�2#���e9�6<�}@��%���b���֦�Hv(�Mw���x��x�^�s�k�Rͣ�{7�(�Ia���A���i'�%w�EƧ��A�D�����^����7:s��үax)D�@i�d�װ_r�3��|�!_M�Wb�F
F;\ M���o��~���N�1�j���$�q���9��(*�Q4؆ݔ����ZQ'
��5�FU�4�������̐廒`*��C�׎��V��$��G�Y�P�n|(�r�i ȍ���K�	�a	�oT)��iݓ��uts$��^��U~�����g̱��R�d#b�⭳�I�i�?fDp埗X����o�pF{ل�NH����v���(	Q�2kVZ-��~>'����5g����P�I/�h�m���~�f����������Au��*67�����Ve����/�Zu�,�SJ΀����R^����fʐ$����l��Ǯz��c��`�G��n��(�y�E�舨t�=Ù}8�J�u_�_��2��
��b�\�[��%\�-Qr>��D�_қX��&��Y�Rg;C��u�+��f��G���}8���M���z2ܺ7S����8'��H�7H �4~N,���Yh0w���k���ʖ� �o�h%?6�v�5�q��z� d�~|�?�����"R���)	��"F��J=����m{���k�\-X��*ե�;�>����c�z3�za��F���X��\�q�~9IJ%�f�P�� ���4i�7g����*w���)�xx�εӅ�G�4����N���?��S� ������tIE��_C���H4qHc���Ǉ #>wVQ�(��4@��2������>�
�bk�
/�~���ms�7%�|S�V�k����� u��x���SL�%���:�қ���z�{�*v�cT��0��x��H�Y C����叔qk�by��Q�`���/%da�1��.ݟKn��C���^g��Ai�����4�^h�)��UXU�"NX�Yb�X�(� nQ�R#���x���fc��j�/�Y�n!��H&%����������NpB�p�����e��r\<Ο�\s��"�|P08]{���-;��}�&^]����+�&I3�6�,��\��� �����gCs�6��53E�	�˫��\^b+�����(��b������҉���j�dý�����F��p�c�qM�{¿���wK���Ӯ�����z	����v&�<�R��͢�c�BW��a�W�>hI���U�O���Ğ��E�"���+W�9Z;�o|�;H�{r�
�(һ�1`s��J��c�A�룕9�?`\J�s=VAAQ���gN�'���g~��\�Ĺ�J����0�z���D�����A�1�����|��`4<�t���*�]���i�,{t���31u-;HyI���k]ӂ*gW�����N��ṟ9��'�Y��������zф'Uڗ/g˭�@[̸���>ފm�hp�V>��7K�#�9ʫ_���s$��*�}$�����ևG7Ք���)z�2���z?�ﻃw48iP����@�( ������N��1W��g8hH�	&@�e˓��x��R`*-z;|rOZ�bP%������H�UX���xy���*��A:��6������Y�=T	�J9��b
3�!Q�Y$��c8D�jÖ
Cw��B~�^����J����6�庂�.��$��g���S�1R1������xZ7���h�"�!ًN��	�7�*?���]%�P�����≊�1G���[�յ5x����o�%��T�H�t��yЛ�Ph�{pt�=��������3~��b+W}�uFH��JE��}��SH��.˨�����x�݋I&�Ԡ�{.�H���?�Ĝ�3`|s������V���%�ߝ��y����G>?�t{��ש��ܺ�a�f���d�)*bN�l�JK��j�AJ%���!�;��+��Ptƾ�Cp�s#٦Tޘ$���pk��oC�1 �Z%R��3�f4pM�6�%	}ܢA�ǔ��%��Yb�mHC�O)�A}�F�o�Hb���P��39=F��V�
x�L��#���}]Ǳ�[tC8Iz;��xI=�87�ɔCʬ��R�w��A$�z_������ �{-���8�.�I�tk۸G�g�'��dܺ�*e%)���X���t�{�:��n��I�E�Ɨ��*9$� �����J��]�)�V�|٪��d�J������S�)3��c�V��CQ�zhw����l~��?tK�`�m���5�Do<����,�sZ��c횋����"88���ݒ���wE�C�7��ډJ�p�P�-K�c˧��E5�Y-�R��N��<�\���CEL���^���,5�Or�d)[��K�KE�av�ҏ��#|�A����ކ2�>p��8o������>����ҡ~�r!T��+����IM����{OŔ��F�QEt��Md��і�M����wq'��b��φ��0PW��"��I�h�t-���#�ަ���T��2�?�_Y�A	6��3-(��.�� ��'���x�6��5���TI�$�^Pޤ7y3lW��o�X�/�J�4�nb�`���c��V�g�gt�\�Zov�!�}(`PK�n��j����xV�Lq:����X=�g��f�imh��jG�7{���������S�:��2�����y"��n��jۡa@+�YL��ș�"�M���Y-%����C*��D�k�nv�-������ql���g�ܚ�m��_��+^QP��0�FA嶘�#(��OL������=w"�{�%���L�n��PdaښT�6'D������V��}YZ�)T1Nr2a"���|��*p�@_�]P�J|w��Na\��OG/�L&��t��&�A�����!�]�u��c�t�5ydw�5�����6هX�y�1��������*���y�%��w«;IyW��E�xB�$!��R~̣��\̫�h���>d�R,h���Xݧ��6(�f#����P��]�7�k���믎�pe�-�b6�"m5̾�ŵ��|@�<D6��/��.�z��]�a����)�r�)�9j�Vn�_ۺ$-��谦�1AM�T�kt�Z߹j��N�~�����x�45���.h��� �2Q8T����cr�#o����ʸ�6X�`T���$zX2�r���Ms�n����H�����OU0n/D���J��y�1�v��J�٥�������{�r(�f���FY�n_��!���˭��p�"���	�qh2�:�j�R���v%�˦^�����V��#�T24�(w�t�J�:�"��HX�)<�t�$��fo�W7q���V��a�9��E'2�yzgԲ=��������~��X�yRb�k�����wy��,x#���^Q=8���g��f���[�X��Q]�!�^?�-���-�H���r���,��DV�r1���[���KmZ�r���|@�ѧY_"]��"����k���X�&F*��}���|�7��4r|-�e��q��_u�uUq��A��d�vp)E�sYaU�>XE�pj9_�TA�OL�3t\M�g�#Q�.��C�wIw���P ��Y��&���@t��=�k����m�5���e]H��A��_-�p���*n�Ů^t��`�Q ��W�Ѽ%�vh�О�:7PεM���J���"��ZOO���i�L�)=qh��]� �g�ʧ�P w������<�\��|��1�͜�V6?��0�RHf�˘}!F��Mc7�s�I*�8n.Mt��M�XJ���<����yR�2�{aC��.W=�'_��zIm���=���OY���^]��P
p��M�[T��	k�ܽ���m����wt���lN��GɽMI����C{���Q-�2e���el�t�"�A�gs�s*/7l{�3?����sW��tL9^c�zIk�n ڧ4bڀ�	����0&%���$�A��M�}=X�A8�"���)>#�����*=��I����LEM>eɰ���&�o��̔�*C��7v�{�"��ePlvɵ��81$lu�OM�+�nK���[�̀��]r�l��G�%�㻂�D����kn�Ɣ�6����VjT%�%
��v�zU�
��A�( {HAݖΤƍ�}�b��u�.������
#0:6���Y�o,֘��)����M����.��L�$w{:,{����U[k�?����� ���� �#�,ݹ���P�/�T�ޚ.�.j8���d��%c�"�y�L����?�{���D������.�j���1�&4�E���Z�k)a�iO���v|���h�D�F5� GG�7]����Ѐ�<��$�k�<���F�8wl��حE�D��X��E�l�{7"v༂s^�٬�=���V��8�1���!�vF<�ůj��GTT��6��PA痫g�7�)�2�o�b�O�4C3� ��q�۩ �4�w�@���F�4�3҈�^�ۖ�(�1���A�P�:b��%��.��-�%�O%���2���'m��>L�fi�M.-��BPx�n�N�������`rB�7����i=%Y-�1!�%tYT`3��S�I�Xa�+�p3�O�Z������.o�
�!.;��st1y|K_O�_�7Ra`\�M���d(@����ߗ7��4��N��8u��M��$z`^!~�b�S@�_za�Ϥ�ɳ�3����ss@���<�$^� ��4�����'���#b�K�f�x�O��醗�k�T @j�ֺ~�	M�q۵ΠO�-&�{������,�fF�w�,u	�6)��U5��bR58WYz�Xői�[l�X�ڔ���,?0���_ڠ=O���qs�$؞^Z�J3X=��ՖW �&'FB�E���
CE���)
?PI�+����a�ru�e8q��0������jnkM��<9|�P�;��q�s=�����B<��3[��kG��``� k�H#�!7c�O)�偝��G��cT��1���4mY��~���!�dJPF���Hm9��0	��|��͇P�^�w����:�U��o7s-�q��8v�I�฀(�s*��W��<�s~��yQ<�s�XԿ�/DP^#f_�"{}�B �3G��@���b5�FN��>���فF��[o���@�^5U�O2Y�7`�:f�1X�u�8l뱖E���O��-6�=�vp�ϓ����Q�;q���?�bI�B�ܳk���J�W�3�]�Uz]����!��6�I>Ķ\0�^M֜e���=?jX��m�/�sE����[/W��l.f�����$U��
����\ At+?p5�v�K�f��]n�\�RH��UY�Q�pZ���4Z�'�@�/!Q~�5�B2���}$���j��C{��Q�M#bT�)8�����>]�� %���K�M5��<�%��k�"��Z�0�C�lh6��V�3k�@������bJ"ȭ�ܿa�^X��q��nD��a�3Bu���eS���/�V`l4{%iY#�-���
Xu�G6X�B$�ݥ��^��pvq�N0A艛[2�_�����=���.> �Lr�A�F��}|�o� 9�ĥ��y�س�?ۗh��ߟ8��m?�Vx�.��Q�4c�B��i����)@����ԟ�����K�WY泿���jb��ڋ�\3c�&�W�w���[�(��YÐo߉��yz����G?�
�2v|��������UC���&��՟�B~�:ȴ!bޓ&+���9 l����̮m5j�i��W��&HCu���]�u��)/�:ǯ�'����X(�G#�8[��������\8 |�˞����? f"�IE]"&k%¹�e����)qQy;Ft`�_��w�f�}C�F/�Հ�2O�uQ6�:������۔#5��FZ �1;�>�O;�"K
�K���Df�\���d�V����Ӏ	���	�3֪�qL��~!4���� �{ܤB�r��%n���">���wz3������e" ���[�!s���Z�U˕Ȅc�}Q�x0�s�4�;��C�T3V+����`P{F:43Dr�W�̃��.)��6	����މ/�5�$���'Z�c�94����l��b|�~FaQ�2a:~G�4�of�՗l67={�� �XG��h8���ٌ���<1�$<�VC�� +�����嘶����罦�T�{J�3��JZ�'�.����{Jl��g��9��?݈�qC���'�?OR ��
 W�\83	 b˩rS�jb���w1�_ʮ���o�e��T7}K��pg��������|����-b`x�^�+q����jiԽp�lFA��dO=��ZG���1�}��4�*��ȴ)f��!�E�3�@z��^L��=�����+�S��Jvq0wS��|��tұ��HC�
_�+�̊����>ĸ2�A��c��2���V^��an���ڡC�.$?�	gF���X7�Ȅ�
\��+5S��VU�ws�zg�6Z�!8�5��m%̗��1�L�~���P6��F20��XAkvJ�x \2�s̓1�˦[��ڟ֜XI���91+�2	|�rE-����p*1=9��2���Tx��a��X��H���?(�1GT? ˦9��fI��������$����`)9���qd���|�t�{�'�>��U��aG%,L�����R�J�ǙG�]��l�y$��H��k�'�3RS�PD���:�3ڪFV����)��u �
j�p��hDW���!�%W�*_�lnZ.a%:�MZ!d���Ỗ�D����{�8� r��A��A�d4�.
t��5ˬ��0�Pka׺�r��R4���>d�y��.y[��Ջ{UC�W � ��Ѣ�c�r��n$���4��fhH��3�i��aGHh,�:yů /�&4#�y0;F��"%�i$0�@Ml���=� ��y�ۻ����g-��RȬC`��Oy��-�:��r(�\8����-�;���4�7q@�:@f���oJ;ȿM��~1�V�����1>��	��c�
�� �ѝ�d�,�Ve�^����>*;�%�<R[%H�v0I%�hA6����)��oz�4��i5%��2���˒����gt.��\�&��Hb��9ېc�!
b�E��ꥺ�Ѿlɴut�E� ��*�ݻW��iZ_�8�o��m�O`�Vf�:G�˙�(���ܠ�H�}���ؖ�I�4x77O�hXmyQ��gU�7�9?���d�$	�~��\B�Y�Ԋ��	n&%1����|$^���gpn-;H�U��9�9�@�4NVu���Bݶ�%˻�.w_J�D��2,�����E���9�}�MN��D�/�7���һ�B)+O��Fn?9w�u�;��	kX�Uh�60�������;���If�.\�D 3���5Gf���=E93]v�t�3''z���؍ltI1���)�օ_�lP�]����r���[�a�U�&w�����IF_�
N#���ufŋ�}`~"� �=�9t�X-�K!M�\Q�AӋ��i9i+�7��	��n&fHɸ�����8he���1��r� /v�����gI�D� ���#H@�g5�8�H�f���I�O����9�&���J���B���I5iQ�6B�`�B~���!�M$#Vҿ�T�GN)`TǔC��6�O��7Ṷ�e��#ck[:�Va��=�M�\�f��f]�%F.�<�5�T�	-���P)�FBK_=�����,LR��>��DjY��:;��[o��+L����u�y?��0�{]o��ia� �V�� ��}/����Y����,Y�7���wx��r��G���S�7A���%�Q����Ŭ��@�/����+���ջ�
�ީAJG�&^`���}ն�ʬ(>�&k�Sq�Ч�ֻ��.��2|������"Jnj��aSXj��Ð_�o+qG~�٨4[�*Luy�BE�][.��1�Sr�����4�]��	��D%t�e8�t������J�@�z9�>m�v�A����ϭ���1؛�$aA#�M��FP3ҧl�����O�d1�|o�Ɲₗ�.FԨ&,C�y�����/� Vl��f-������A�U �8rF��D��,�iA t���b�Bk��L�v��+��(��r�)�$����w�/�X�� G�DsH�,;\�&n�%��!��:�*���>k��E�o��=���G�[�fx�M2a�1���J8���Ԇ$���A�g*GE����������ٕ��ٝ��)�bq�<�H����J`�.��n�� �K�NISd:a��K���a:���Mb��� 1�Sh.��j���\f��t�Q��n�r�O�Nc��̎���U��¦�/�/LйDB�3CE{���V�>G� ����y_Ҧ��x�>�X�� &����O�'l V�?���Ή���0\}�@����Ģ��N(�"Yg�Z��� ���S�.ߑߺ��X[c&�T�B� i����
 .�ǄْG����]����)����(�M	�Ȧ���ɽ����S�Y'5ʽ%a�,�^���f����d|}M���v�t}Ͷ�\<l��X�ٰ�xX�w���7<r�C��m���Ν4�C�ī0��s��`���:�zCt+�J��G�!\��Ȯ������uw�6!N&?��0e<�	�i�ipg�����և�g<� ��4ga���+A�a����-�s�L�k������;�,c��� f$���_-�h҉�}p�)Y�(f*í=^n�ӤOm����1�a��4d�Zk�ӕk��P�/B\���Dś �޿oo�;-��aQ9�k)9����h�u/����\�6�h��~h�QZ�q@���T�_7��x�%�+;�ŭ�՛!H�smV���7_����=����U�)���1�Б�~���6��g�T����r~�C�uh7�uy��y��:7���:x�վ�����`HX�����f��W�!�x����`W��ul*%*{R ���
�4|��n���أ��+������h%��{&���͔���L�7�u:�ʺ���rw|ݜ�^#;�½;�'b`� �yѭ�u�xܵ���r��.�6�7}�'��P]J4E҇����29-9I��p�E1DCAc5�y�������U\�(��Q�p�}�`��ܡn5p~��g��Ors&���Y�F퍨���X)��虳���̛>@�UkL�i��I[`��C�.��O�_�����p%�J�c�nC"3��T���b���k}��K����O��UI���o��T�_�$2���E��ڇ�UA062j�!%�9����œ���[M�_Z�Jyp��F�33i���8���%	X�]-��Nz�(���-�3�r�1Q.A��ZG�s(���Qܺ�U���O��%���C�zB٤���2t�����LZ8..O���S��p_T�,;B������`G�Ӣ ,`�� ����?�3ʮ(����Hb�6��Rz��M���g4��	�h���~�̬�֫<�����T�L"&��+�������.���Rz���_mx����B
��bD&�0�i �;�<�qٰn�ט��֦�����m��F.�X|s!U*�98E:*5�*C�|��: ��>��֎��%R�)�+����S����p�
���~m<�����5Γ���s2#T�7�cX�����?��q&{���C�"�X%�)� ��4��b"�)N>��.ٰE]��#�d�5��)˝��ā}�+���\!�e*��"�sy���;�͸�r�*S��&�e3J+e�&��(�-�����6�^zaHũzT��"����Z_�i&䋽�Em�H*�w*ec1�\3�\��p�}�9���
�����i���`W�Rk����EW��6s��{y!��]�W��7n73�(mޜ���YEu��r��\η ���{�-nCi
�K��[��1�i�/MٰP�>�{5���R{В'�,����rp��we�Iđ��=~�'-H���Y.Mv��}?N�r��.����n��8�Z�q�S���f���8����?(��h���Q��HN*�+m�e�W\&�l��E��N��>�! #��]�N�ܴ It�
p�'.�*�߈��\9	p瓴����1BcP{[+������M�(�iiy�4�XrIF�'���!�B愣$`G�����+d�d���r�� 2$�]ӧ���h�x��%k`��Y���N���@f`��uoa
;DT���K�"��æ}�s� ,6�U�F6,z�׹?��	�ʓ�|�cg�
���'�.�;g~J���^��>�� �"QQ;b�6�ɨ��㈾��xE~gB56K���XJ���:�O2NsPҚ#&U�}]{�[T�I����Y4 Ƒ���it3����D%�$峈��#i^A3)g�lb�d��w��va�BV�r���`��{��l ��^jIG+}��0����)N��I���{~CGUVh57���G�$E��8m�j�������k9T�8���	D��L��I���	|e���˛O��,�hw��y�+�� ��쯦K�����~w�8�5+�Z51Ebl�/Y�R<�z��~8�>�y�&)��5$.o.Ə�:�Ȯ�&��M	�cs���ϝ7�zX%�ݸ��ʘG4
��d9Ք�Ɛ��ib��-��tsg�ĺ�6�+KCe:#�,�i%�߬�S ��������/�rm��M�4Ɉ���l���,+S���}��r�>����Il�>;�&<���*��;
(TG�M��garۣ�w�F���>�	H_�Cz�:��J�z:�&%��~cc�宱:Ϻ�=�n���^���nё<��]d�#ǳ}����#��v����j^���;�U4*�˜�c1�9�('7v�μ��@]&�h���.����u0�Y�8�X!	đT�����ߵ-cH�	R�t��ڵ��p�!�p�P��o��q��d5k
 �X>[=��E;�*?���p2��~ה�IL����V���:U������:��Ȓκ�B_oq4Y����Dͽ����t����q��J�~y��R���?N�k.�{�\^�\�J=�[�����h�0Ҡ�p�u�z�/-�������@��!{�Uvh^�䐖�Jj,=��\��V&��ًvI��е�A�X��5�'�X��ܓ��Ч��º�p�UՐM� �!��
��˖�8�
[g&1 t�ֲ������B+6I_, ����2��{O��,H'mi_Z��Bw����J|p��<
X�Xu�&��� Ӯ��j�֢;˯��x2���X\�=;��>J��]�^��֜���<�0�>/a�Ak}-:Hq���Jl� H�a�-�cyp�BW�7�=��M�QC&����²p[�ʹ�]J-?ёbptzq��X��	11�  �r�z��8�x�$kb���b;�2N�6T����$fQ��`��r��r2�H�|����9�Or(���c��F��ug遛�D2��GC��'LAp��L�q����C�v�T����X��'�'�U�o���,�ș���G��}�[���Ɣ�B�B���t�%���E���H���������W��%��\���&E�X��k��V��})4Ǒ����U�Wa�"K��6U]�b�*�0;�����}(��ش�gۨR2���C����p�-ߌ�qו�tf�mr`�G{�զ�"m�}r���Y��]�
,�4ܦ��Oѕ@3�3�a�r��\:�{�k��I��H;EQP�!�����ߖh6:WbW�x�� :��%���}�I�q+�9�[��m~��@���~�~�Ǣ�$/�ʩ!C��szQ �J_� ��[�tx�	
.��	r�Y�K�)b��&��Խ��ù0�7��4=�Ev	%b�~4G�(��o���F.��i�8��'�+P��P��:��4������^���}Y�8%nr�g�'�.�>� �ڜ� ����'�f��xXen��\��{C<�	K�I�+GR���l|��8A�[n"��7�3Z����x�08�)����E{A���8�a?���? G�tT׫�>��(�u\��[�lG=��p�5���d7*6�KR�=y_s�U��'ʞqny��N=�W��~��.]���*�O7Y�����c��#��G�q�+�슣!H+�K�[���/�bvI>t�p�.d��r(�5�5���F��B1R[25�<0H��1�QCqEp�2�`�dg:Kq5���N�����8 ̸v�5Uoc�m���5_�c�!���=<jh�T�6b�����<�-�$w��\�T�i������	��?�ɋՖ�#l���k���m8̦�O>Q$�e�*���q�]p�n�.��˷Q�����%�=&�g�`��L��X
8�&_M�9
֠^�>���b�"��P��iq��4[l��e4�𫈣��[B���3I]$���gs
�e�6%4��
��ҢexF�a"��������������,G����e������I��`�[{�)�d#׉���C������t�g-<�Q�����U�b�G�S�e��]�e.��B���M����.Ӥv��k���6g��X�CEvl��8<%�Ð�z�螥	[Nt��Xտ(��G�?r��w
�asl- A�<YiT�<���܁7�fs�a8췜; �a�Z����Wo#S�KU��z�?���,_>���/j⵭�*P����{��-@�~���|����D�j±����4醝��l~I��lG�a�e��2a��*8Tq��m���J0����|�q4����4�>Q�ݠ9ђlYf�!��/�^��ƈ�?�����`iY2z"�m[6?v$p~� ��P�^������G�8	QZ�^���R��ߓ���CE�};ܨ��Lm�[]%J�,YÔ����ӕ��uFרo��U1�N���x�sI47��{L�'�K������+��Y�nÞ���If�H�8�<i�X.C��(;�$1q�Ś8b�U�j��=�l�������S�l���f�	�A��ރ%&�}*�n�e�.ˬ�W��á�S��`i[?�e��J$��ˉ�m؍Kc�1o��P�2�(#�G1p�)�k��h�o�>T���B0+�w��D��P{�5��)'��V��.�5�'�����d>�c���ldz�7qme�� A���^S�O��I���'�X�����L=��.����˳%UP#����D��L����[�Sw���h\�	~'!@q.��)o�5�����k%�R���K���s�aR�NA��%]�$��G���h�θ�޾rH-#���B��Dg�;ԛ�~�g���2�󧑜����g����f>E5t�m��
��3�/ƕ=+�	,}��r3�~�:@8�H�	���b�^;�/�u����k�8��_�;��ޗ�ƽo��N2�������)�����T?�7~oW|�.Mh�L��`
0� �u�����J��܋�9!�~˂'��SMߵ�+L@̍+&�����R5�b듀���H"ŧ����j1Т�6�A�{�<"+K](41�!.^/��99�>�a���bln��1@���3H�k:��Sj{3��'#�:�D�b��P#�	��i����@:3�	�6�^�CS+\e���)ǳ t`�1��l���.�p���cZ;-)�0��\���l��k+��R��Q)[n�Q�t9Q<9AD|�F�@���L�iWe3n���� ��+�%0q�z��술�Gh���`N���?(ٿ�s�p0}̢rB�<��,&���H�h�iF��>�>��Au9�jT�b\���������W~M9z�T��xS��U|1FY��qRps�6��8C<�9��G0��hz�M޹F����0(F���CI��5����E
���K�S�k9y�����Otp8���A@�󇉿�H��)�[I�VD�JKԫ�R�v|/8�3r�Kg�"ҍhS��E���DĘ7W���NB7\hȤ��uI��I;j��n�r�6�߶�u����=tF�����k$��t�#*v�~��`ˆhՑz���X��8���68<���ѿ:p-��M~6ݏ_��hdm��	��U?�;�cv��v��\���/)]خ�y����rO�&o���;+��A�71���~�,��(S���֐�ͤuF�ΰZ�
j�%��/�{`���w�]ﶛ���8�o��nce�!�"�!�d�~nE�� ���^8�=5��n�mB�W���$Ƞ�'�a���9��R�!���C�g#��<nͩ��<��5YO���J��|A�N%q
���L�����g�}�Xo��������o�`��0M��_��#�I6��C�"\�u����ټ,Lh��g��=�������7ǒ�-��$�\3Ѧ;����� 4�7��/w���Y��8H.��d�C]�VMF<w�W�C��-#9ߊ|W=P,H�*�;EW?�B���$��'�I��R�Dϳל��lx9����b�H��R����&��N�,���߷0�r/<o}�nv�CHy��Ȁ��b���)�J�p=���QvZ^x.7 ዘ	��b8�Ǒ[ ����_��?	��a4�L�C�>.0 T6�M�c��8��AysQJ{��6bч�[��6������[��G��������pq��AT�y������Lѿ��G)�1���+��� ���r���^U���l�n���y��yC!�eraэ/�1�Ȳ[4�� ec�	�q����tF�7F8�yβ0�����S���M��]�F�$u��Y}�����?
�����匘i�i���$r�w�k=�G���"*���
�b�8���-Z�a!j��Wq�ʈ�՘�'�/Ԟщ5BA�������%<x�,he�Ep�c^K��:����GN���JXZ{����'�����Ɯ���.(`8�`�9<�Mo����|���c��YT�A|�UnB���]yK�K��1Z�dڐ(	���[��d��e����c�n�iR�ˢ�Ej�D,���6��y�7�_@g���I��v����R����|��8՞a�ƥ�=��S[|� ��bȂ6�0'9�����k�6�$ �d��t�X౔̠|��m?Ϫ$j�TlE�C�/!a�i�Ժ`�K;;N��L�b�T�f��ݟ��)�]&o���5�!�A���E�՛Vg���:r�M�� �����5.�w�,v>��@X�/^KoJ�H���@�������Xs\c�S�Do����d��b�M1,W�,�O�T��a�7EV���꧸�p�ka�֕u6�	���FR�Q��cP�I �b�:�tp��"D���tE�;X�{ҩwq�1T��k����u��h}E>3
��f����u,l��ߟ+�s̂���D��w�ɂn�����W&���������{D���$���!������lW�
�Q���!6�W�}`}Py�t5�T]��F���RRо����J�H>�A �]a����pn�ҙ� ^	�c�����?��b�r�B��	G��l�,b���{��n���S����l��
�Ǌ��%�8�����F�*)��Q�����Bl��6�K�m͹���p�1�:��}��n�ƺ�����[�Wn���
t���xS�^�l���(wK����l���Ay:���|fR�P��j�3zF�#	Y��W��Yߌ�	Vh"`z��=��<�w�K,��.���h�]dȌ�2U����!��yI�ٛ�卯�h��8��q#�e�jo��o¾J�A���a�����@;�j��ڜ)�:i����#F�̄�5DR�+�g+�7�e<�U��ڮ;��\�/aC)��K�V�-V�_h>VK>���rU�6��-����q bV��d�2�s2ZܳzA5)f���L7Z��^䉅��}�лH��LP����՗-��'����@5�8�E�>v%���Gd��P~���V��o�E�>Ԕ�8x�뜵}���ۃ�ٺ:"�hz�'�8�uY>�G4YC	������!*��L��DֆY���-J�C����d}���1�V��遘��li����9���meR��)��́���6���c��KEh���ة�{~O�|���E�Z�b ��I$��%���dgr�.�ױG���X\��V�,��i�z��c���+�t��=�	u@���4��{E��%��A���姹�� �
��FE�6�"����{�q(Ej �c��o�&���J}:�;d'+_�@5/2r]pj%�r�ta)3?d�`�^W�GK͇ў�����r|Rd�\ȡ@؆�+�Y�pY	��|��K�d�K63��_NV����\�8\������L_~BT�`�P�����;��I��l�
9*,5	�=nϢ���� w�+r%vQmo���!d��a��-��	�!_]ǛF���k"��TV�v�ȭ%�M�$k�|��KJ<(+h�H���b�tep�¼�7Ŝ����PBƒC���ЦD�K%�;�#��U�O�ҳH��寊���S�do� `������y�8D2 �C�8J�_j�O��8F��mcx�`���`�*׀�X�b���*Z�K����jN��������x�D�ѭ�Iɓc�2�
&X�����x�>n����\��L�ŧG��>#)��g�1����Z�|O9�s�8��%Y-�W����f�d)Ǯn
m#��4d@��Ĉ�a
I�0�A�t��B��D���yd�Y!�cq��8#GlO�ݱu����uP���4S �B�����V1˘Z{N��i��9����ݣO���ve�bEC������ʩO����zj�=s3:�4���5���V��gTV�e��\��d�&�U.|����]=aPc'Y��c��*Z�������0'G�-n�B����a���P��J�a�Y�N^p,(��%�Xr��^���t<�[#���N�M��R���t:I���}�����ߩ�s�h����%�)(B)��,8=/Xn�ˁ�iC(�-:��@��NZ��8l�Ћ����GUR}ғ�4�V캲�JA��w������Y�N!�=iq��">]��z�����n���G���6�[��e�ޒ��a����-n|[n7�\�����f�� �����B�TCu\���.�q0�h� ��zlS]r�'1���qB�,�;�zh�{٢t��v���J!ߒ'���=q%�_��qVt?!~�^i�IC�2+%m�A �oMwX<>�nkj�xk̬ڟ��*YW�wޖx���<��W�t��K��)�6�0���P�@LT���Pċ��Y�~R�L���9�`4�cܗ^k��R�t*Y3�J˴�gԧ���+���SSj	.�Ld�~+�}񮶴�N��i�ك���M�H��o�t����h'S��=e<�~"~W�m��g�atJX�&.@EKU��Z��hG��ލ�����n{��3��&X�Qt���[��k�F~����,�$�	��i���ŭb�Ӱ�G���c� �#�T�͇�Q����4(d�a���z�4 �!�#0Oq�'�~��"��B})A�5�ȖU��E�v��Ɣ��\7�k����w�#�]&w����O���
��@���^��?��[i�'lb����a^��r N��(�8����µ�)y���7���\N����I���^y!םaQ��ǀ� �U4檕��)���c���w%�'s�&����˛�[��J�}Ki�����1�G��A�k҃�KEPq!��~37ѩ���r��ә�&��{�<���|�D'G��@�9��m�";A� ���H�E�kr����q(��0(��}z����:$k��
�j�td5����hkEĂ^Gt@���a2�i2-hj��+ӷ|u��0k��d4<T[��䖟Bf��g���&�\%��6^4�B�z)l�J�rkӡ�7�=U ��$U����-�x��v��?��d'a��s] �?�Y^�Kq��t���J� H�*j����[oC�{95�]CW��B�Q�볏}��9��<������Q���W �o�Z��C��t�c�{��?�� ���3�-R�!	q9���qU�ӡ _
j�9Nؚ&º3:���MS�k�Y��;zKT6(����u�'d� /�E�%�+Q��o�i�����9���0E<ɵu�<�r��5U�����r�/� ^Jܳ�;:#���w���G��ڦ�C�\r��&�wń�<��Jݜ[��5 �L���>R^@�k(�1�` ҹ�:�3:E	TȮԤV��{��)#�p��8��{�:���8h��<2a�n}L�x��L�<��K�r ��C��`y~�v����i�H�螸R7��X��p45�?+Xh�3�˯��D瘞�kW�\�*��=�� W�1��L�	��c����Dȁ"��z��EO���.�3A��B�R��yq)�c!�{f&����7H�_��w���B��Ca��ͬ`��D)�4�iVj|ذ�ݫ<H>,ic�d�Ͼ�w������>��{��!�0k>nM�q���3���'������Vp�أT��g�:�`������hL�hrX�[S��I�R�[@��B7��k6>)�[l~w����2V��l�_���U���%_'�T�g����k��^���w�c�H��z�`���^8�h����D���W��+�'9
l��=쓽0�s��i��0�rگ��a���읻�h/5����w��^���Z<.	l�Ǣ��ɝ��HFV�;idcf��i#���mQ���:�mF��zw�:��I�v_�-4����<~uˋ]��L��!���V�ï_*2)5[����'�Ŧ�3E|6`�U�9�x�>|R�{����M_rfצ5���ǝ�e�����&�N�;�ֽC�D�3���&|���3�� ������UT�m����F�WI�.��mv4��f @\���Di�n�A�&gH:`�6ZT絘"L��h����cp�Q�T���0{R�� ٛmbv���lk3��D|����1�G��)�����^����K�n෸����4u)����Yr�,�!�[L�$����q��*4ll�
�e)��}��ւ�T��:`�ƛ��������-�l�M��_IbN��T���.�h�nj�b�n:O5@��	�	i1x�;V�!0�_�̧�+��xx���d�V��9J���F��W�8?���E8�:{с:�^z��BM�DBd�/א����)�,=�W�mn���łR���;Uધ'mM�M�B�Ӽj�v���bX<�(t�B����P�DG�g|7�L�'���

1�-yyJ���r��1,|i�C���,ݑ<�}�޻��L�������ϴ��zP����h�����,�B�����N/������5�ϱ�B��v�A	�:�Ġ�u5�KcC>��뭌�R��<��Di���=4�t��}�:u8�R�;f��n��YY��2<;��-$W�I�ܟ?1��-�ʼ->�=����ݱvŧ��FHf��]�ز��<x���ïv�'>�2��G���I�t��^�Ӥ��b.��������C��^�"�?�N���MM�j�?<۰�4�k���މE���Պ��1����;��ִ�F��x��֝�W�34��+�N�:b��oo��m�z��7�����HF��9�v&�1���.Ry��dR���S��I��$*�ߜi���;�k{�!����Va�_o��$O)����e��B�\(�]|�8��{׻(�TExF�JIw���r��1w�Ē���;0$c������Q�%ob"Z� oP��F�a2�I��z��k�^�|ōz0y��n귙�dt�� �3Gc�2���˶�?�k�Ț�������`揢u4�������XtS/�V�Tg�g%xoN�:u�|���Gp�;;��ր��%E�
��gU�p�<0�l�9a.\|��N{7�y�O�<r�x
71a�O��Y�W���|���E*M;�|�5��{���n6$QU�����&��p�L2����{)E�k��Z.��~�ѵ��� ��n[иʯƟ��Ѭ7ًt񓝉�#W�����B�w-Ճ�o�!/�n����@z�f�(�Z�l��t�T����Xj�'PO�֓�Xl�|�3�)��9-h�v�t�)��u�`���@F(�{욅��E�7��q��k�3���G-�{9��b��#e��N�� ��E�A���Ԟޘ����ˇ9���nv�������vj������DV���yפ;V3��TZ�}�>�f(�?�Z�ދ��2e�mN]�����&�u����Ow��D Op�z����!+w1�������H�Tz�ۚ�?\���� �ϗ[�sY�q5v���na]�<a]2P{�t��m�ߏw�+�w	�O�ӔC�j�?}n�Rj�,0[�m��F�����A�F��lqE%b�wT��1-rMZ�s����=�6?}��/O�ڕ}��{���qz�{l,��:��.�
�pK�K�Pq܍�;������N�tˡ�)���;�A�6[���iV�����9J��͢�q�3�I.��u�Ke�uG�Ȃl�%�U՛>h��p֍,:��u��Q�Mʈ��j�YY�ɾЋq�h��:�e�����}~�z?˜ �h]Ϛ]���ē�3�0X��	&��gp�rW�'Yx~Ld3�F�@��>m��c��Y��{_����l�����x7���7�''E+��S��t=>����~E�2��}�8�\��		�iB�Fk��$��g�4W�Ev���%������ZMFVa�cje�&�V����Uv�W/�ڪYh���P�y��( ]�)��U+��eԸ�^���4[H5钗�x���Z̝�L|��IɸĤ]�m*"�m]�g�+�R�� �t�7^p�#e��Qۺ8�2i�$9�m��\�n�N�<2�������6�&�{�|����D6�]��+�r��A��"#�ENӈ�]��ͦ�����?m�
~v���st�p���6׭����7����th}��n��9:�#��C-�}�����Y��۝3�������x��Dq�k>I�W�,o�5��N�r��ض�ɰ��O�a��%e:�	��:~�8R��JԾ��$H��:S�5���tL�gM��ɛ=�)X�vjF��L!Ȇ1B#\9}�"��V�բ�9�B%	�Lj��#�'�k��?�B�QH7&`/��Xt�TBж�o�Ud4Ŀ����`��.�	ȟc���f{}3i>���B�hFYi`��Įya?��yGvY�� �IT\"��+�~��^��+���n�&��EK�21�6�An��9f�>�}��>N��Me�\5���\U�KuY?�*^� ��SC�vc�����t�P�[}�GJ��a7�It�l����u�_5��L�9��Q��۶�+��=�pjZ��X�c�~ƴI]����N,��b�`<&U��u�Q�[yay����@Sg2�ًyu�p�ٺG��.��%[y�u#s���V�+��M�R2��V��yc؊p��-�t��h��75�x[�MSA�Ea��e�W?@:aQ�}���hNmctl>{�؊@<��@}�B�Pvg�zٯv��!�mچ��T,0����-�U�V���h�j�`i)��o��eX��ʣ]��rcd� .u����&OB�xp�D�m>�#�w<�r	դ��jiK����hh޾��0������!
F��+\HB��$����q��o�v��e��\��L��@ݫq�SX�1||����oϑ�o��K
�Kw9��D(E��b�2C�:��H�
Yle��R��S&^-Loo�(�'X(�E�2��BI���х���ADg�OC5JU�݋D$q*���suan&Rh!�D�*AA���T��Ő(L�a�e���s�b��ɀF	{vW{�^M��jSu�qŧ<K�
�#|g�<*$C�A��0k���7�~
,�+)Hg6����~y��;��'��5��Ѷ>ʋ� ֳ>��{1}vrau����2	s���G��HWi�J.�@NLzF�3�LFW\]W�+cw��Kuc4���H�t�P��?��xf&����!�+
Y"�;�[2�q���C���_v�=��Z���2m�fRx9�}"YC�&���~k�]6�ҫ2C2��Jm�ˬ�ֺ���Ϳ�s@(��,ي"U1@�%�HKK��K|��ś�P�������m�V��e�!��o^�|�{}B�l�'�4��)wtP7.`����EN������W���5آߠ|4�O9���b��pu9�xF�����P�޶��V?�,��F(��6!?���D��}����W��2r� ���|!^��?|����Fb���f�	y���k�e�J4��������pYD�XU ��[��*/��'|1�k�� y��������\	J6$��<�ʗ���L���<�OT�d��v,lڍ	�weO�=)��Mm�R�#�KUs+�i>U�� �K}���ߠ�*߆R-�(g �{]��5�R\/�������4F�zI�� �u��O�����6����%���қ(�+��ݪ���X��o��2Zq�,�������PE�R��Z�4$;������� +���I�	T��&�����[RZtݡ��Qޖ6���T�.�L���`�˗�oz�ꯦ��h+��L/�8T�Z�R�l���y�[2c��H���uL�7�����JF��L��8�ϼ"�1�7�4�{��r��
�7M����p�ɹ�e�ֲ�"%N#@�t���5�~�b�Y]�Q�ټ_����rE:��m+�ز��鐼�ɲ��4�3�1�EW���E&/ѯ>_��R	֤׳J�Ho�>��B=?���TX�F��\������[�L������L=�|�Y^stYEł$QA@��.}D>���Ӣ�����D�d�9��f{A�~�˽<��E��1��Ɉ�:�k��J��񦻭�'��o# L4��Ɩ�3�0)W�@���QȆ�C"��P� S.
!�-��O&��N�]���a�yx^n��Tڕ�Ԉ���<��BL>K�yNjq�c��r�����"L��p�g�!�5�<Fٜr8�D�h4����%�˭�M!Іax
<7����4��ō��y��;:Y����iF�{��e6��\Gރ�l��9�M,�gt�qN>�Sw*CнB<
��NTL�v���n��VJ��F~�7���ز��Z<�F��(��Y�
���.�~Q�j��8DT���GOPU�	f�wa��8���Be�_�][�b����{	�n��f8���Y��_]	A�n=�ؔ�ͯ��%M)��*�9�r����t���FM̞ݐ��$J���+�4-:2�4�/�a�l.��h{��4>B�@�;+[Į�QJ'�#��s��#�$�8��.>�����QB������\�.K������>���u�}����_�흾d���fv��ď�j�?��5 �%t.Н��[:�I��bq0��@�tCl8�y}�
z��ӂ�t:{�S��@�D� ^�~�䕹$5�N�����=�s�����V�v��~�|�bE��;���z�Z8m�?!�i7	��Q�[}�[��{
R�,�9�{S��p�� ���	�>]4�t��4}�E����Ra��_1	�z,��̘P�hz�zT+������������1g0�n#����6�Q39��O�.��؉�1r& -�l��ؽ� X��Va�R���֡��8��i�I�S a�w�w�^ZT'ԽM�4iؗV=u��'-ڛ$�����sZ�`jc�mxilۧra�'rMs(F�@��ѹ�T�Eiۚj������-�${��G�C����l�FMl��Ȣ1�-�/vAʂִ8���`��
��5��ލ�hֆ;6�:��(��LK���c��SF��WD�5���X�B5w��1q�cT�"�ka^֡U��HTdh��3�������11���A.}?�;�,���҆}����y��EuMW����'{��=�d�'���+YU@c��>��}ѷ�s�<�#�⺄���s� �R�m'-�!��y�򵊬�GQ�k���ǭaC���^��q�+�B�
T����^�,��5�>�A���c��ȫ
#�k��{��'��|Y
�Y�q�Xu���'��Od �$t��/����,O
&S�=��^��Y8	�		<�wcP�7�!��]˙p1�⎪x��|ɄqY��%3 Y��9��T
�|K	26|��+��-W5%��ݍ��~2$=c���?z�.����Tvi�e�LCU�M���BzB����G��e�k�B���ġY�j�v��6?x;��q� ]��T��T=�p䋄��:^Ps
P2����>��7����	�t��y���>�;�5���mF�5=1�ߏ��OF��YƍY�]��h��_���Aѡ˫=rL�wB
zԜ��M#1���>���Ul�L�^�/�S�	Q�hZ}��	J@L�Ǘ(�0%��mN���k*�"�&=�ws��ZTh��{$���E�o6�lN��P¨wnQ�q���c�*'q�=�
����v�m��[�3����M�p�L�h� |�qЧ�R{�Ul@�~�)�=n���ˋ��E0\}����5uP}r@��eU�?�c,������x��T	�1`+XdO��f���8r��/������_Ck�����Ff�F)��R+��pҕL��EЏ�$"���ׇ9ὼ�R�����F�io�(>u)��چ��v�R.�H�
˂�k��b�����w�>�g���q��ۘ֞��e�g�rSD��B�'ʻ��P� �g�4�P��(���5�Ձi!cvqU�"��0�L�^��)ǩ_�k'FbL��B,'E�
1��L��_MI;��1&����cG��G��x�)�ט
�9��&fZ�a�N��E��.�!�)k���J��sʤ�6�K:N��L̩¦��I]9j���w���W:��q��҄���$���#�aY�7l�+m,bWmX6���S�4��=.�P>��xI��{��~O��GC�)0�+�Mu<�A�9;X���)P��i��A!M�1b�89P�B��%�Y��F���,��p%�F���(S����di�?
G	�:�(���#�������Ї�1{xl$��h�����-F�v���^w<�"��ʧ^ZC8�aC���_D�'@	t�����n1���MB��5^�oj�:�X>�L�p� vҺ�^���D��}T�B��`�U���=��`� 5�GX��B�4�� ���2����>Ԧ�m�����t�C���:�Uo�iBgWѡ7��N�q&��xfU~TJKEڳ}]L�?��) �=Y�Q�/"E��$�/�t@���G��&�2�(Cz�8�^,���9�)���w�1��
��0��U����p��:�==|&�x��e�F�C�")�F`�u}�\ u��Y)�	%L�ٴ���e0�8�Wx|߰*M53�R�1R��,|���ȧF��q�n>w�֪TQ|)x5�z.i�'i��D8iу���:�(}6�r^g��}͊�<��d�q+#R?*�fDw0h�0�&ޖbΨZ��v�p�NRZYw���C�[���
��m���M眊�1Ht`�Af� �[<�1K��g��e1h!�fc�Y��3ʊ���$]7S�? ��\������^���A�O�W�F�3#��Oh��tV�*�g��O����
���׽x��%��b�Hց���mr]�����������< 9�~��Onv���[i�mBU��;m'T~�?�yC�1���0�ֻ��s~Q��,k��ݵ�^�n�	o����Y(p�S8Jт�z����d���PYg��3r��c4���1�/��r �j�m���i�(8���?��n�b��5
����	$nOk"Jn_�C������m[�iO����B�a�M��+�d�w�67�c���&/��QxS*���g�d�͎`�r�fa��[ƻ���~I�D�Ti!�,{���.���!(=U���'N�V*rI2��kQ~���� ��7-,Α!<c�e�1���ǽ�-�h��;90^��EQY�0�
�
�����r:{y����n*�`�d�W{V�n��bN.��tiz��>l7���/��B�0�|��؊�l@����6��6]އ��'ʉ�@��Q�����a�}��Z��vvb�F�����3E��d��F^_+�S��ӏ`�} ���3��&�lH���R$���t'�w�U�X��[��c��a�1��e�dD�D��˚�9J�.	�s^�_���KB��<� �v�kV�u� Z�����we��5�L����J�](���ͧՔ`���]�-Wr%�W_�㵷��Ί2FH��.k�2��U��(�Z*�w'�&=='���P�^L����|ϸ?f=����������L����mVKm,���2���uwa��u���p,_�J�'~R)�l,�,YSY�"@�v������g��'�j���`���Ag�I�"�B�oNʓ�ΛZG#���(�sEd~��K��L���B�td}�������)Ym-�tl��="(���ȈP�~�	�  ��}�0��_m�]�BpA��T�'��[ꝋ�������(]�p�	�g�w��r�MpJM]��-Q��'�
m�ZS���XC2��3���Ӵ��w�pM��gU��
=�g�ߪ�6�<��,0/�,�AZe��Sܿ_��w���nN
Bv�>�φ�}��oE	i_M	�~���9�f��U�1����p3���VɞN��Ȼ�k|��cx�/���>����*�"�&�s�j�&�ܦ��u5u=�7��ejeN?�Q��/�&6�&{�ۊ�� l5g�W~.3&7�X�(�����\�vN�޾R�:
����\�޽��u��7��H%��F
�H��oi,���� z���fVa�}��P������B�<�N��a���X�̔�,��0<�������wS�b9���ˇ�ǛKv�/L�x���S.Z�}�g>���T}8"�f�]to�XL1�?�)_O1<L*$ўr�w�C���m��8�o^)�ĠX��;��f ���e۴���\@&RaS����~�䜩�IC�n�4�E��b���b �͋|C�5��>����N�ku)���S�G,�t��Y�:��_���]�)q�?xC�E��w���-�ш��Z$�En#���+���k��+�̼�k����t5�F�������q�}.s��WV�`#���
�YHr	t�mk�%���ӟ�6Cc,��g�(�'�Wϔ���B	`0i�9�c��e݁*�3�\��V���*�Ī��b4��`<��;�DU��l�P���b�r� �L��v��n�f^��S���>hv#�������n��q4Z�w;C%���;W���8�Z;���8��;�c4��Ey|���H?�fF�ľkm�<r�������u]�u$)�D)�����C=]a�D�Zz��7R���L� �V�^����o��fo-j���Ǩ2��u���e��.�1�K�w[W��D��#�̴j-��t�%*Dꅆ�ݡ�<�� ך
��a�=�F�Od������S.Y�'瀲? ��R���w9����������7IOށz�0�fq~���~�m�(kF��=����\��,���~�,5.;�猿Baa�R(�u�2���lѢ����#K3P���]4�~|�Q�1� �X��@e#,���~��[~��c����Y��$�P�MƩ��}؍��à��UI�>ܩ����Vɵ4��c`!��.x� ���|��LԹ��k>�]\�YE�n��$S�H���)��׎D�`=96���<�oG?]���C��HT��O �+�����FN�y ?��$�v���{4�F��X�4��+�����{�Btoo"O(�}Ÿ" �=[�4��fb��(��6�B��ǅc87����k77`r@�a�?�B\r_�g�xc�զ��;@㥔�#�� y�N�÷[)F��گ0��a��G�^���e=΀��s��41�$H47=��M�WϧDo�=�E���������`����My���Z'x�����	�!�T
I��M���YF$�����7�s����fO���S\PJ���#�'Ǩ)�W��ڛ�L9k�·`����zz���*?�B@�E��k��1`.6�A\�i[�71��e�Έ� %��U� U^T���)
fghZ�f�+���Mn���:��7]�n��n��H�?,k�L,���c��h�Z�eAЮJ����jIgc��"_�_Ĳ7+�� �NR��7<�k��ڄ �8l�H�^�+��LN�1g��<QK�NzP4&t�����'�F�����=o�v�p����s��-�����4�AA�QA�T�g7���?���9s Wf���Q�rޞ|h��@�͉>%�c�`��Ɖev��PG����<�2r:=�<j)���	�Ȧ�����_��Io���0��c���H���!B� ���*l��aM�ô���������ޗ�6l�ٱh��F0�RK���g���&�,�n��	���E��2��dU�");�4�~	0�l��ae�9�y��/wt5��+b��r�9QИW�J��_RBn���Ē�vC$9d'ys	o{KT�<������p��`�7�?�g'E�e����,�U�_{���ֆ$(�"B�0�{�-�'do�S��ѵS��3�ˢ��\�s�T
9���.m0�>II����I!��M0�������"���v[�2�����<g�7L���Ԃ�f�ɵ>��3y�����V	)��|֜�m}Q��U��I����K��uA\��V�}p�6!Z,2��7���0U�fotiqjU�t�TE	�m����h<Y�:�+�))��'͕&�+�&�Ğ�^	�{3��X�V`�F��Y6��Ś�<�A��BB�
+�0X����{�pJ)D��qoD��c���D*)�1���ɦ�m˩�,v���ևj�z�B��x��M�97ـ|��4	#�R���T�7"�mQ3>�>5@֮���wY'�fc+e����d�P���/������<^?I�-��"�O�Π�3;`u��b��^/e��^�4" `���4�!ϗof2�e<�?���ܧ$8��۳D5$Bn�[������#u��r~:=�UU��L�J�N��If� ��3���L�t؄�,��E�����i�=#�����H9S�I��YX�A���5xau�L��������j=7��s�rD~���!>�_�c4F�0BHѲ�1���5.c�0k�)�~Ue!D�R�f kʳ�3pVC�����d� ���Z���8:��N1x5'~�K�#���w��� 8��;��Tg/@�> ����ҭ���+g!K�������-�G���]o]�Z�'�"M��ۙu:6x4��p��-È��]���V��F�D |� N^��ïD�������\�u_�M�aw�p���Bs�X�� ��|�C���RA-1Jsɂ�R����ȷ��O��J�;�?���`����x���+FG7���ͧ���A�*����j�GԱ��ա+%�ͬ�l|��$��p�F��k�P���5�t��ڰI�R�����2����=�E�]�U�VAh>:+���*7o��P�tz��<��
�l5,Z��m/6���Z%��Y�៭�g�w�O�i|+���귫?�䈂}���s�/o��׼�����̀M}`ƚ����R �0�����jbk��_td��4���yz��I���<��pX7��*k빈&'�n�QӴ������i��-�:<� ���`���U[�"�kz�ŉ����=t�ϻ^�)ar=�<��"v!c�G~�ȞBYD����"Z�;����@R8��o���.3?��$Gqwqp�e[8���5;US�%��8r�,~�T_�8���R'��c��>U�!���#��Fغ�T|q��M�c���ڠE3�@D���~"}�Oz��.E��(����)���u+!\ `}�)hoX�7�#x��ئ}����Gt��3:n���m�ׂ4�[��7Ay2�g����iv48_p�/[{C��Z���1y+�����ʯ����^~�4�:�!�|&g�Z�$���0��=a�A�%�H�pU<_�F0���z*���������,[E�����k['��!;> ��Z45��3kB���l����`��"ud@h��Jv��[������N�7=Y�8�ޖ���fUl�����,�j�M��1B9�3#�	F��n�K�\���	��@��"��޶L�(�g0|
Մ��[e[���)K��Yh�vR��l��\�H��j��!d��W�"�����"�C�|����~�P�F�?���^'�r�Y|�2���P=�r���eƷqV���J�<χð=ҐGO���E�y���q��/ti:�ߛ�oB?;�	��ZY��=h%��`&�I>�����]���<U�4U2ʕ������Wq�d��g#��Hf�M��K-�8�޼��֘������'��$����|1���wuuk���p	� ��v�����{n����v�X�H�M��(�oY0<�U/B�~sK�?��ʏgv ���!J��͏_��S�QI|�a�'�F�K�|�a��*jd�v�� ��d�6$�=؀im����?��v�{|[G)�k���	�y!Hj&��8P�u�m퉄�Ɯ���χ�ɥt��a9�����d����p�t/�Z*���DlT�8�|@ި�!�6u����=�|��2-�à�*�{�BO�bd[��`~�t��-���f}^gB�C_
�/��~�GBu����/�m%4+Q���,��w���܆aq?z�=��;���&�.xd�`b)tۻ��2�P�����_�M�}o za7������
�K,Pl���a`�p��/�Ǧ�Ic��WI�8�I���s���������0����M녀VɃu��B�c�2�fa/�eU͕�L�|�'I$��y��̪�x=I0��w��	���I�W�f�P�F��nKպ+�˫j.��T�djT�F�O5s��d�6���8�<`����dihd���U���9GEs�z����O&����W�k]]&v������Ю��_ؔO����`}��Xn3��n�����{4� >Q�r�j�HɎ�l���;Kw��vC����|P\)@H�ݖ�yխ�A����O���WtB-ӵ��P
L�	�Dn��R�,rT��t���9
�xIb����ȿ)�LOt1�,�]lzZ`����@fڜL�J!D.�ȱ�ʒ��y��i�h;��{�k�Nt�׍@b�i*��U�����72�Z��>R�J ��� ���ǋ�	*.Nݑ�
=y ;){e���C � \���@��-�c���]���?J�A�\��|Z�5���hy����]� p�B����3Y2հ������:�9�ڙ<��^�H�xW�5A��P��_$x��<0��)�cQe��I���!)�'�D	�֫L(�E����Z#E�����a�.B�i�@
xw8K�x�i�6'����O�,Y-���T�	i/�}[z)�yT��:q�<Q�ap�I�섀�8i��G���{�e��%v%JE9�ك��U&�EǏ��L����P��%�&Nh��\�ʣ!כ��'��-�v�H� &;���l�$)��J7A0����$�@/����t�:b�ͪB�'��#�6Őr���4�{�h �|�+GqmO��.$�|r�D��^0��e��N�u�0��f�R�?�E#�&N���I��{=����Q���kحn��;���#-��(E{��N�a�W�֦'��0�mN^��ԍ�
Uk��/2�QD����A�~��<T��m�l��!�K=�@��Wj�ONS��9#�l�(�5�bb�v4m�����$֓W&K��o�ӄL�!�d��|�!�mb{!�A����F��W6�V�f�q��fed���T��@�#��B��O�azL�Wi%^��R�]Q��� }��xry"S��^Xu��ꦋDVtv�P�\VEg���ew�l�*�h�p
�y,�\ ��8��3`;R����|a&�� <��ؓ<�ų��E{U�$�~�h�7?y�̆��c�J��	���g�v_��W��L-+#H)��$: �@���x;d%�e���]s%���L�j'*�Y)�e�*����ҥ��+	J�#*愘Q_�
�Q��c�8��4������wh��U�1���7 �y���:����t[���D��G϶.a��x9�du�h&\��lpu���n~��!������Բ����W<�T9��f�^ԖP�o���q�
��ƺx���^����G�3��d6(�Q�ьr��.�5O�5k#睢#˜��W6I`�oLM1i��]+R E��d`hj��!��h�9wm�p���@��"�d�.͟tNq��æ�G�ʅ�����~<�����F�7!q:�ti���։\�&���&Ш�h�T�)W�Vz�W�v?�FP��`��i�`\���A�h��B��M1Mq�<G�"��	�O�J�����&qh���c�@�UM:TD�e���0S�=U�>�`8���)��"�\vU�ڦΑX��љ7�zѦti�~�J�����Ƽ
4q���#c�(fZ��c%�6�A[���D��͂���3�X�26X��&�E{�^y�BKS]Nl%i��|b�iFZl����3ہ;�?i���*��'�𿝀Ci��TR��S��b^l�}{��-�c�	s�	R��Sxf��Lڥ�ւ�3��NK�pW^�ֳ�Ԟzzb,*�ӿ�:ѡy�Kj�Y8q^p#-�t Cu�eȧ�g�|q1{�/��}�[�[2���~�F8�<*��N=pDP�}�Q{��\�p�Z����Pz�7qT?6~5&���V��M�������Q�0�^4��4AVSfѰU��%�9��at�7����� ��}9/�b_)�����ǴgsedV��[pݨ'������۳��G/ݞ����5'8�4؍Î����ۦ�p���"��&n�[�n-��"TS��
e�*�|J���h��E~#��3��2s?��x��Ym�	�ӄE��:��`hM��:�Y����X�mIv��R�#.��)�F��u0ҎC	~ԕ9�U��jI�O~u�-�>��8��x�1�$1�3W����9�Q�Ӈ����E�/��Z<Ҽ̟�`�����^Q���A��I>�!N8k)c���NaJ�ؠ�ђ0<���S���}�ԿJ��wd.2���+���.�K� 0kvd�7ƬgH��9۵-%�y0���s��٬�k���4�N�4�Y�^|��^H��h�"�4�'$G�����2��v�$�?���])<�֜E���5:ߔ�N��˒'մC���u Ƴ��Īa�rDk)��[>Dk�Y�	�7d�P��\ ��x��E�G���a���߫�8��=�+��$����2��ɢ=%�)���1O@�=�y�#L����@O��A�ݭE����$r����]L<�9�1Ey��&GB�*}��Y>T���P6٩�#_��͐�����f��fv L�M�+��%��,Z��x~a��4�.*88���A
��KѲ��G�6��U\ԟЉl�7mI�t�x�]bg�������$��ܟ$ ��m�_�^]I����5Y�������,Zᾭ)�����P( ɰQ��uL-!Qi+���W"]��'Rd��-����o�?�ёK۹ xP��ި���]V�0��4-�8�F�������:��X�����$�t�t�j�ME��h���{t�i���EƑ 5ҏ^rsKܨ��Ƈ�}:�Ȭ�8��@�� �ۑP�wI��}��v.�o<Js�?�\���9���w�5Ɋ��K�b�A٤����ϡ�Y�XG����^�6;��Pv��ts�r 
��e�\�
_KfM@S�3G�%���湹�c�d��s\�8ֆ/)8.	�pEt�:Ddn�1��{�,	s�͸�!P��	\�U�1~��yk��w�fr,�/�쩌�ْ+Y��P������*���Z�w��s��� �j��M��
�al����E§KG+H�M[�7e��d(?�m���4	�������=:jW��9��а��H�{���Q��l5��!��cX��0�JC|�f�Fn� E�1�!�c�[���,��ж��o�	1y6|&fe��W�C�`l��f�tkP�C�Cs��l���ko���d��"�[IwR>
q�]ea]��
��M/ټ�Y'���u1���H)ŎT�n����ׇ1��NqCo������g�a����E3"�"�Ia�s���P�r�M$�窟_x��P�'�Kl��*'��0�9����-'��P��/�hf����Q�3z��{7�zz3
��44��>�r.,�"5�}��j�<_��8�ժ>��<x�@�v�h?@" ���&SU]��r���@7A��=t�Dvs��a���@	��v��=V=]^�����j� �C����3�[��K��[2��f����M�5�}Owsl��><�nʜR�Q��r�`<�c�(����bUZ��r����8����q-qCW���W�7@p�ʺ��c����9d?KJ�V'�Z�!�4 Pv !�5��6��t��]�7����<<g|�8^������?�Y�@7o"�K,g��^��r�L�����V�?��l�L�fӹce�YR�<�Q���pCw���֠7A�.�G���(>Uŵ(�<�jۃj���Z�d����ʊ�����-W�,o��>o���<mv!Pﴗ&�m��`��=a��6o�g�C-�P���_����`�-ⒸN+��/��C��lr��J�:�ZY��$V� ��,�	M��}��R�ƌ��jd�?����y���﫬���/"�(D�~ ��W�h��|DF�{e�n�7i���w�#���?�u>����9��ì����;��5�g���)4f�)�Cu��Ce�E���M��y�����~>����r-�D��t����M��5mj�����mr1� {G陴e̊�+�t;�$�h��&���,�G=�Waa �@q���O$]p�ۀ��.���v�Z�gg 7ԯ��x�������k�0�&�N�!�^����CM[�ȓ��<O��ԥ�Xj�`�T')E��9�@oP#�T���O}��v2�B����R�R<΄kO1Jq��G[�و/in1�8g�g=t�������d��|���D���[:_^�.4+N��ҝ>����-{�R��"�@�Aviw�T^ p[�MT�Z��$	d4�n(�oń��r��6##W�)H{��b�A}�GD��ǩ�⟶_��TT~��4/��S�@_<19A&��_�h��1ag�����/8�0JD���-�^`u1�[j՟��1�հ��)k���y���y���Ѱ,$���q4G�t�vN�6"��[ń��s���Ko����W~�T�I}p�O�%�U��� W@����,���2��"x���QM���k�Ic4��c�T6l�]�v�����z�\��y�Q�)i�;����6����'�>��_��?y��G6ot4m릴Qώ������TY	�*�wPa�vl����_�0���F�.�����ˡ��7��O�a����k���(��)�ü����x,��˯֐R�ô��3�#�G�:��JX�c�7ۚ��D�pAq��h�����c���5��~�1�?�р�Q�ߋ����l>�m�jq�󟙲�|�4��L7�hMt����Z&�4*-?LJB��\�y9�2�N+�S=���pjG7�X����KϠ��v��;t�#8��zA���¼���)�&|�B0Gօf��uQ�%F|EsD�ƻ�9!ă�l�>d>,L6�>�%���C�|�A��M�7F2�\y+B��+�Ōv�2TS�v�R��>)ŵ��~�"�x �Q~��8tD��
��e�v6Ӣ�[8��H;�V��^<m�֦�@��/��-.:'�"W}��K$��c̕�:i�Wp�K�K�%��jY.|CY��~��}8�	�U�e����Y=׬O>^'����B���`�#\>���2w15# 1�A�;�F
���T��(Z�<�sB�rr���ey;5�k |\��|4�U��>��EW��Z��=�/��1<#_.sG��?��)�c^6v�@���&�s3z7��	��1U��^��s�/]�Ձ�~��E��r��'ȗ�[�a
7��#���AD�w�V ����2 �<��j���j��ѳ��<-��OUcc�/�kM�}��a�t
�a@�ڦ���:T�ʥ���z�r�����h�� �` ���4�v�!�Ar�nlP�qF�k�ʨ����0�83�E��¤z������P������J�I��@e�˷�ʼ{��l��h����t�8F��
��s��v��T��?�QN�˴Zdz?QE~|�1����m S���C�����W�<��*��I��}-�����=8'.���s?}��:_�?����Z�=a������%��
yZ���cv��Z2��%�8?*>@c��L�/��r`��Emʶ�!%�){�z�kHC��1V^������"���\� ��R�f{Kg��,�����[��c+��4H����]�L���� {��#�~_���v=>�Q�-O�J��S�]��t��W�����;�z����F0��S��_����JJ$j1,�f_!�)�I�bK��D)od��4��Nn��R�b��bهY/fJ�h��!�w�೏��t�U��K��t��R%b���A9���ʡ�J��˘:(/��0�df����!P-2��=}v���a;j�I/
j�2st�8�tS����t%LЛ�FR���dO%�v׃4�CΞ�Q`�nV�+��`#](k��ӱ�LpVI$�߭�.�YU�9�wkU�?��q�0�+%7\�5�ߡ�~����5�\��|t�J�����3�0�J���𡑲��8���Tݑ��\c��L�]�o���:�3�{��e���6�S��,��3� h��U�7�]���f�q7M��;%���c�2�C׃����2^�r&�V�]�;�ݵV򖵦�frX�X�vv�՗�t�l=tx<�<R�a�(UŇal*���
� �`Pg�o�Ct�����JY�&�V������-тj���:�@k�Pw���R��_��31mȄa;��&9�x}$���e�+l!$�Ӝ~��U���8��Qj9n*�0�]*)���B:��K� d�Q��B�]*�XZ��b�L���C�P�V��N���r~�E1����ͧ; �v��a�O$��[ Kײ1�%���P��� t_�=itC�^�㘔�1� +.�.�a��f5.�k{�E�D�ܻ=�+o�X>~�6�{}>�G�;�=�4�4�l������4�&e�B��m����5�C@;�(<0�X�'i�=��H�Q��+��#��aci��aq�	^��CGq�f�"#.@�X�6d�񀽀�N��ׄFwe�En3����N\��3)�������x*�Y���?+��4����ڐ��4��tq�l�����}.�?��Ç�/�������bO�P�f�T��lX� ����D��ݞ5���=���Fkf;7꓋����`���[�ŏH��62{_V!2f�|(�����,:���B�~�?�	E�!nu��ih�#Ndq���E�]��e�YМ]Ut
�C/��Pj���x��n���д�k�A�m�O�m������ηM�`,�axX�〘N�pv�
��B�	��Ex5�I/x��*����D�t�I|����W����`q��y���zF|�PoJ��i�ASJ��Kz�DxP�K$�09��9x]�v���&�>
��] ��o�X�M+ޅ�]��;?;B��C��0 ��D��WM�XĚ�j�D�ށdLe��F����A� �5��� ���w@G_� �m�/�����2|5���JJ���ʈ��p6�F~PS�]��/VT���5�,X�����������i���鬻\�06t��j� �V�d��a/� �c�zI�x�W�*��y2��w�T=��s>�0��%ۺ�܅�'Y�Q�fu.}[T��p���ϒ
&��.5 ��/+��\[P=�_$�c��4�;8/�.�B;�#"c���y���5*��ͳ��������+��c3������1����_�����=8� �tY����5_n����ݎ��Z�1�`�C-�p�S;"l%�����n�1ә�풍��o��������H�[F.��什
���c�#l�����I<�3�[�5U_�Fh�1<W7��79#;H��@�<h��;�X��h9������5�|�_��l%56�<�:�1��tz=�J-�U���;o1�Zi)BfBY�`r���E�ޓ�{�=�z�/�a�$�>-("���Ƿ�,$)r�|N��`o�I!�'���G�vk	h�|ղ`��[{D���ٱZ0���V=͍B��i��\��ėj�*���5奅�]J8g���SCj�Cxb�06�t�Z�):��/y]i�l��(O^��K5�����_b.�.��Uѹp�����H���|�I���.�ŭ �)5݃��\����k(���~�xh�q߃���8x6���q���*�	�����)�}a% WEN����yB~zb����!bw5I��$P�+�|,�>����${��]o�!?�� ��"]�/Ǉ ȓbݓ�M̰'�{����,Ek��A\zՕ��
W������M���2�j�T��=�֖u��Ē��v7/M$X��/��B?�r[XO��������B�{/'K�����K1�������º��cz ���foi-������4�0Yk�dy���a�ݎ�	P�욃�w�!�*�3:)�c�0����H�?ҩ���@����S�#⚇��f�3?.&˭�F�7 ����C7(�����k���V#��bۗ��%��ߧ�m)S��_l��K`ՠ5������]�����,���l������)e�N氎g�D1�b Pjݘ��
���l�ILOe�^lx��w��ƚ���nh��!Q�i�G�5�>�����
6��WGf=��)�m[/:j��т�**(�-PH^��t>���E/����2�!��m���l�f8���,
n�CZ+I�����`���swk��T����r������2H�	���g�q1a�B&=�&�za��k��&��sͪ�b������aw�8%�뫜a����f�r��n��DRsl鍱1�=��t�[B2'�(�tE=֝_]�h�6+[�ml���}|/k�X*e�v�iZ�	�s�o�_��vHɧ���8Џ	k�C=$'�	� 9a��3.XZ6wN+�H�����υ��`�bMp%�qs�zE'S�Ԥ�rZ`>9�7Lێ
�jR�*��q�%�����*��jD�f?I}���
ļ9�dҡEja�*��d�F���ƣ��7>��h�x>�cq��.����]����It������Z������(nUK	6\��վ;A]	h�xU����S�D�oݎˀXvEu_gh���'��d��)����G�E$)��GvA��(9ݶm=��2��SEb(��e˺vʙ��`|��w+.�{�NKyw�o�b�Pv��ԍS�j��C}�p]�]�F$&�N�b��C�e�����Z���g{r
(X�@�Y�J6x��&��,�=��
�92�]�ZwW�Y!�W�eۢ�WM�R��g�ߨ��������ٕL�/#�b�s@AŔk@��vۯ'A�ʴ3�W�3.1�I4BGZPN��ऄ֔�e5������U7O>ЁLm8UL��v$�����BY�f2��O�us\=��q�-���"����Ō�m[�!��o�3|�iN��O��#L��p~ x�G1�3�c���2��v����9�!�~��9��6҅���M�'&nHr�Z!b���"^_6SP�8e౞A51���X���˱��'=�8Q� \�D-�I(�`PV��s�ip&�*$��O���!�O��7�'��#G��P<y� /$H�R�u��knAk��)�D��
J�87F҃M��]�i5��'���񊏚y�	irz�,j��[!�M�]WZ��a�lǂ��h� ��WR���!oa��%��Ъ&%7�?�Iĉ'�r�qf�� ����_�_]��t�楟m\�HP���	�UTx�����q.?I��I��;�����T �?Q��"��Z�Q�o�8R���7v�2w�@�^��B�S�0�_�Xeg?�[�<$����|$�Bb%<zC^ӊ�:�o\���8���z=j��8_����X����V�����rF�ʵ�c/���E�Iw�{=��	R�օ/i�Շ��!�o��Aq���g"�������(1��IxhX�h:� ��Ypg�N�g�|sB�{�2��$�ab�b�����y������i�h.+�;�!I�=ʅ�f:7�5.;ք՚~��F�Ѩ�Л�$��^�bR�f�2��Li h�֏�v�H��Ԛt{����v�Vd���F�wɆ�����D��	R��NQV��i?���Ff/�I)P�O͇!���{�HI�l��g�Y�;�� oӹ��9t���Iگ,�f�2��޺ò8�*�\W\��{y�M�S\���G����g"G<�\��CvEb���_���벁e�c�.<��`NX��l���Wy�^�p������ٳ�Q��zA�P�kDX��Jո'i|�9�[6�f�*I��z����T�[U�d��f�;�bk�JݐS۰d���a47���c��x�X���V�W$ g���_�R%���0<��
H���Lʭ����;���&��Tv8�)]�	Jє{S!�:-�o�`��W���@�b-6�}螇����>�`�\�)�@��j.o(j��܄vb�H�n�� ��3��Yx鉶>I�{�+���Y�k��3O�u���I7��6ۼ?s*�o3F��}���8ZC@��B���y�<P�i�dsh�$�����΂P��E��֩7�ZE}�3:J:�9̮��׼���Dč�jҒs�&&d�C�T{3^��P��%��,Fڊ XȆ�E'V�����c�L|�r#-���q���z�w�ы;�,83Ml`��غS��U���X�Q�1(A�D�,vײ�-8`uS�h����hbNF��-�f��e�З*m����
3��������b<��s�,6$��f�MS<��̗�ϱ���o�]�9�q;U	�Z����V� s��&�{�B�5�O�����/ #��/Q#��[N[����m�e��ߪ��F��ٜ&��]���T{sf %��c�	}�m�O��Bm��!P}
v�H�:5\ƚ���~�h>�6��p���_㾯�}�j����V��� �)�hŚyh릾؀F�Aը�ْ���p�՗��H#:d���Vr��\dg⫻@[ϧ�^��$_��	Ϝ�j	K҉�sY�m�\�q���ƶJ�
�����@�X����o���n:�8[嚐�Վq��ג+A���6�˱�D����8;G��i!u�.Nw������{����ir"d�H#/�c䆁u`"����ޣm�j��b����a*VsU)��bm�����p�t�&NU6{���8#�$��Y@�q���^�QT�=d^7`�ɔp���\�h���SI�Eu�R`{v\u�6�}_���>�~`�X�c�Y�4ϧ�_[5���ND+����4��
�0,Oa���7��߷� �c�	��:�(�I��m��F � ���Sεmu�
"{���q
[9)o*���v�%ݣD��-��k�s�C�,N���=�^����+�۾C�~�|��B���iAQ����_�����[����:�z[)�91�R2�����PÊ�z��`�<���s���rM�C��ٳ�� �$<��j�ߒ�%��X��_k#d�{���>$'���	=�a58���<h��*&��n��x�l"�j�T�m����{�._��7��m>��I��&1�}��y-�)�W�(b�a!u!��-�[&)%1�����X�N\l��ƀ8"%���ŧ-57��A@� Uf��t���xp� ���v�lh��	��}?{�:�e�������'�rE��rp�X��%=�{h����@���_����т��p"�&��ur?=0]��ީ�w�䅝����x���{����k�)m��!�Hvٙv)�?����ЉZ�q�/v I�U�q� O���ج�4�eC:`��A?F���ԙU�:���	Q���w�2-j�M#�I�j�s��Q����=Ҹ���L��ό�ZH��+t!�8���x��K��($����L������&�����1\`�'��^�׼�$�5�b�E���ro�2c%�צG��>�랰�);�g�4A�ZQ���}��J(�6f���F07v�\e3ZH3��>@>�3���W�M�ཾw�m0��@
��4c���|���z[���U���]��A7�.ꏙL�����N3�?�ڬ�O�����[p� ���ȠȏHZj���]̧�Q#|R�S�C�b��C����јB�w!ّ~:)/�M�-���@x��0"D�2X������EyQ��7L�s��+���ў>�����0��!/: �]{�Z�mI�o(�i;aY�4{�W%h�� �dAR���H噑��U�0\d���3�7m-k���QSv>;s^7��c]4;�\?Lu�P���+����T�����k𙁓���G� �;�P�0�lrx,��@��ג}����� G��wV6�`�0���^��G�N���_��k�̡��N����YtHյߕ'��$�踂��xÐa����TU�mk	tR�{�0�@*�3��� ��+wv���d
���[��d�$/�ü�L��^��U�Y�F�6��阦�!'\�j�1Ԋ!�����*S�`����͈^�w�f�l���J�%�9��e~�T�S�b��+8ư�ׄ�SjB4�u���{S�������!n}�����E�l=�k0JR�X�	;�<��� ���������|V�����8��<PɠAV���Vk���}x���m5���jZ�fҌ����r�ݡ�����!��=l�ݔ�ޤ��r�ߒ���Ʃ��<eBS�ֽ�W~�oW����
���Ww���ơgP�:|�iJ7�85�>�T�Nv��T�����/DX��Ų��ܻ�r�b�x_�
�����(ޡ+��i3��_}
nJ-d'��$FvG F�ęP��n�8�r[�T�������ɰ���S����g.�ceݏ�G��3�2u#?�$�AQ���!A]Zt�}�l���#��Վ�CU��9���
G�n�|��	j��k ���1d򕏧d��*�/��J�G��(5�D����G!v��;� �	�k,���O|h�2���x���w�\{����mN��"bl�`�P]4�i~�>S@���|�1���N��#F�`$($;O4l��pѬ����Nmx��
[�4�2��1W5��!T�� ��T�:�����>x<�FŋߘV���ʾR@U���KQ��AS?��R~��bs�	*R6-Y0�9�?F���Ծ����	0vSU2P��6����S�e0p6�!� \2(gt� Y%����F��� <����D[����(��������f�Կ>|��-�� ����26VZ�8Nw�YK�is�A��c��_��wƜ㑺���i��'i8E�Ն�l�����A<29pN�C�Al/����5�{p/&��*�f��(2H�f��ӈ�a��O]F��^�&"��!kZ�t�oM^%�=���A����r����d�To2
�S�r��s=��l7ɉ1L���
)� h�� �Hj�����g�]��4!zk�O�D�0�ݶTx����bN,�V�9�p�b�	�7h�^�5E���e\h(���.b5D=ӜX06p�
*��Nx(��s��ztJF��f��`���ڏr�!��YT_�,NL�������~�P�;���J��#�.��Z3Ǣ��k&�����`����A�WH3���Ԑ�=x���k(G_.��p��I^��m��Ʈ�����������k��FE%5��/?�����{��DN��* ۽���Å�qG�6����zf�&�=�h���ܽ�C��>��,�f����� ��Z������"S\�v�6!��ύ�`�0՞�zk�!^	s[�د��pY$��Q���gE�F(�G���s,�t6%o�iD
U�=�/\�c���ns~e���ںGi��� �,0Vň�Bb/4�ok9 ��&�K�D�n��[.���8 \�>�.����d�olY����Q�Xzb���N"5�K[��I�˘S��z�&�'�^0_,c��r�^=����8�j�Ru�-��n!�X�m(���w1�fƜ6ڿ�io�:�;BW��f���;Z���%��e�&�i�+=*C��s(8�S�b}#To���a|}���YQ�p���*z1�< oO��5�7َ������XF�	�E�Lh�W�,��H6t�?����Vx�&��5H/��R���W����2�}���D������.��������D���;�:����~V�22�K�;��W3�6:S�#`o�)�51��y���H�B�}��S�Rl���$٢}(�x)`���ҳT�]q�ı0W�C@���hg��Ӛ���'o�W�|2��d��J���:V�p��6�(���m��~Z�Q -�J���šʘ=b1�(y��>�;�#nD 1��@,W�+0�\�p�J�\�Ԯ�*�y��/��˶�7�t=.�L�xV�~���ܐ��P= �Y+�b�Y��(��O[bS�2�1�=��X��� ?ayY�p'��`�D�k��)α��Fj?d�20<��*å���{���'{� �ٻ��6�)�3����)�6�$���t�οr�K�6 j�މi��|��Shz����+�ۼLЇH�9�]Q���G��Ѻ寂8"g%\iY8��+p\2����>��T�jѤ���_��˒�8��k�}s�rI0ѐ����Hl9�	��R{z�$�_$�� y_iX7��Q�e��
t��Ǒ�yx�=��ҫ��4oku�Ϗ��2y�j��1���um)���߆y2��ܺ��x�ْG���3_/,�!�w{��A8�8��������.������Ŋ���$�0pd��6����)F����{4�f��(�����J���nݯ�\�n'�Cn��*�2H&�m�G�Si��M���.~R�l�:��L,O7q�p
��ß��-��FOv��5%�Q\q4�B�W(9c���es]e���&9+m�z<�-6�R�쎍���h���-Nk�8ÁO�6��oz6���a/V��㲳�U4)����U��@W"K,U}FW`ꇱ�ҽ�b2��+��s�Ҥ��Ƈ��7�+t.�w"��ݥ��A�6��.SZ�\2j�ڡ;>7](���:��z�-8gS���f��S��'��p�6LE��0�bΫ�r
v�#������(h�O�T얘��v/5�|8��/IA@x��G�\o�N�e��V,׵����"�\O'vl"��Y8g��/�h5���t�~��W���۲�P�P:W��~���P���B���m1Ȣ(��[���I�%ߢ�vE��0��<$8����ݑ�jT'��5����0�5\.Ȝ��5�_���<�P��ڗM���,�+j'���`���ڝTn�`�]��t�J�����}u������u#��w�6(�A�AeV\�\S�:ڲ�.�����hXF�����_��r\����Yh+nM�|���+��;���	h�#|����2�3�(��V�>&�r�xy+@�ٔ��rH��xZS��]�|�G̆e֗�n�n��S��S������qW�4���D���2(uJ͟�جk�hʠ�r>��hL`9���B�3On�����V�$�sVá/�ee0UjV���k;j��Q�4cľb~?�T��{�6j�����;_|(iY��	���PcX����{��~���Ue/�|��#��� ?���jXOb�%%uH1LjC�˹I�t�x��}^Z*���Jj���R('km���j�����aݑ���!d|rN�����LB�
'��6�1��/�'��j~e�k��"�V4�ӽ��	Г{� �N��]�;a\�qb��@	d2U��!04I���	R��QR(����+|�QQ���^�<�dЛ4p����Vt��~B�X	��L�p�0Y��^?ĕ�e�������U:K�!��3��;{��BT<i��g�d=v\��*�^יI &jC|��U��r�*�b��+�"��/��z��6�8�����$�WՑ-����$"�z�5��> w�삞�r0eݙ3���I௶'n��7w~�<��@�SN��՞b#a~��i��%�1��y�+��۬K��7�I�4=m�:x��O����+�]7�a�f���sku8����j{$Cw_�!��L;��|����<>�Z�l�}m�T&#V��6�W�G+r�����A���K�H��r���RԀ#��5YTFO����-h�If��O"cնP�)[	1�	U�TY��8��g���̏�CsȞ��048�=��J� �Q���2����8I�#q ��ظI���y���q2��&s�G�O]�/g}��A���S��#�?E�7�`oz��g;72�v!���\����5=�Vȼ�����-/;��(���@�<�����SԺ���N`�wK���Ee(F�I��m8��B��l	�[�휥$'�K�K�u7Yŗ��V��DZ��f��4�-����D��k��&su�!�}R��7 �u�9�c���u2R,���6������*��j�o�¡�T��Y�T�ɳM=�,4�ޏ��}��'Xa�.�!֋^����j�P�Y�Uއ�]�V>d*�>:�m�c.�\*�]��y��r���@����r�#�E8di�1ᮖ�n�d��b����P�^�ɫ|�����{�_ޑ��(~��x�����K3�� �~=�t����)���/Z�lf�u:�kV3�nE����_����:��!o��z�tY�B׼ȉ�B�����=e��B�������ak�%�޶�ƈJ��1g�Ĉs��C�{�
`�٭���r�x֊+A�ZVχ2ܥv:�⢰�Y���'Q��Y�X=L�����k˂i"\������XE�/��m	�`1d�K��❭��ذ�eY9Ў�)+K���6�Q�fA�y�x���3Q��2��@��A���%ն��`+5*w�s��	��-ʋطJ�
�]i!�P�|��e��r"�lќ���=�R?U�>Hu�zE���mp<��g�r�2p[*8jٿRx�>�FP܎������h�/�r%�Z�{�X�[�y|OU���0̑��e�
� ��!����E�`�����S/�:�GdNAF˻����r���Np����6���w�c0׊�qA �b*w��9A�$,��2�rhhP�6�'��7r���|�vhg<Q���=`+�|奠3���=�)Q��	p�[͢HsH%��w���c"���#� �!�X����0�s%Ixn�3v��Y3�[z�T�uU�H�m[�<T_G���5�K�
��';Tu	�<R,z�!�Hx^��1v5H��C���z<0�]�����,!�s1ǌH��n�Zv��ҵ�(��E��$�hÑN�G��;F6�Y����$��	q�&�e��s�=a��*�.�d��3T X{��EX�D��q��<�bc�
$I�o?�F��3���"p9�}���D�#��})�O�������LM���� r�?�1t���#ee�9��A��=J��$�2V��6��@,vg�|���L���:ڨ��F��y�ais�1��Dz�hs�W�����yjC\{<s��2��4�eQ"�_�F<ڗ�\��b��6�[��H��8*Us?lnS.X�
l�T�7&:�]��}�.@B�h'c|���\�*n��p]/sa-�yߙâ6�W_:����W$�R9�����9�ڒ�/��x6n�
�5/$*�&��=��.�CZg�
/c[���<qg1D��R�?\W;�j6���F�jZj	�ZHrrAq<����h�����W���zp��VK�O�����e�0y��P5_e�W�`����{���qJ1�*k��d��ֹѹ��tz4�^*ZF\�3��.!�����-_Y���dv���7u]�f9%'g�����O�ݩA��&A�.���9 ��r(7�| �BWC����da�>E�F��^�Kֈa���i��/F����a�]	�y��$�;E4n�ѱ�������� �f��0
G7�2|������#@Ff�v�A����!�����P�E�Wa6�j|U�h�iI��=!�HH�I�jSq���Kg�y'wd�������m��r0Uq��	c<��f,Q^��FFr�^�\�T+��/��KE�|k���P��* �0��nW��E�����9K�n�M@�>T�jE��уxg����Ce,/5��<&X���5�D� ��NS8����hX�n��� u� "9���b�ؽ(~=��7���δQ�D�3T�B���ϛ΍ʽq9����f��I�i����]0}��gƕ�{bp���_��Cn�E�v�D�/т���4D��.L�����s�zp�.k���>�M��,�Ԉ�%�M�܎�
�r3vCV����[� 5 �Ի0��h��,��W���e�?�0�I6�0_}A#��}a7�J�+o�
F+���F�[� �{�S�L��bsz�3\�N|��'����+Q�
�y�B�j���R��%G��HT�U��XPQ@�+#Յ�~�F&0��(`�!�`s� ��xі�,����Y\�*Z��Uv�C����S� �`-�)��t/�$�ز�=\����i�!>zH!�P�������%��yI3��;Z�.OAѯ��M�� ��*DiS�}�T�1/ɨ@A8���d��2�<�f��.|1�܆��!O�5��?E�[�ۺ�/!S����71�W��ϲb3�l!x������!��7L�嵍�P�`Y]������G�f��/Ud�_�D�d���ZC��rd���rg����+a�j�|�G �6�Q�P�@�<%�[�ڀ)ү�`܏?W��(4�16��q�b��V���.�L�yJ��N�L�z�ĩ�����mJā�J�4�Ux���W=ߧ��x�Z�^|��=ڬԻ��vG���Dh��Y�+ŧre�U)�YH�箙k�EC��ݴ.�s�go��i�:�K����Ǯ�ܸ��^�\��,�������R�>�yId_�iq(	��t�7�x	�7i�;�G�J���n�}ѥ�p�����S�5!GL��k?ƚ\�N�����h�;�����NԖ��9��L8Lqeo}l�E��_�|�������s���DdҼ������i��dT�L)�7�����`\��1��Y�gTz�v*K��LX?�j���z���[	/j�@w2�@0<��=��9ԑJg���E-��O�g)�Ģٚ��d��'�`\�D�'��3x�mG�/���ώY�A#d�!U�\���Ga����A�����{����	��;�sS-ٕ�M
��|������3�IIn�J���s� :;.`�,� �Ei7��b��<�������L�7��7K�;��"�/u�T���DE&f?@��#7��_	 ���2��10�ʞ�8-�"k���9��6��G�{��d��K������ۧ�����\��x�R��� �$���jBWkh��9��Q;�lw�T�vz'2f[�����P6�O��+���O���sr��ı����
6c���ns��	���������CD�=�����Q��Z��Qqd^�߱D|�Ì �N�X�G�輔�>��d���W���p[o��؍�	\4������m���xa�ٜ��3>m�dp�5�&CYq��HG�`p���0�R�Dm�4������}e���ŏBUri�m�S�a��=�f1�E��Mf!���5M0ڽ�<ma,^��-C�}�*ײ8��fʑ������/H29��҆�/� �Ģ�w9����O�~����d��kn���x���;"�����p�ݶ���u�},�K����
�B���wkq%.5��%�	9��Rh��M��	@m<	��g���p�G���etI��k��I�p��N�'xP��W��co�WX���E��)U��eNe�B�p�n���.�0&�~o��z��|�eP��#>{د~7�?�v��K�d!4{m#b�H����=ɇ�Ǚ�
`��1��r�)rP	fK���N �{��Jú���5}��>����a�}�pb6+9���j]��'?$ �j����U|wn�6ع���#1�nt�|A�p�{,9B�o�Zl��
c���������m\�'��`���yԝ���/K���+⟡�+n�[�d����5����?�"O � ��R��ꋅb�֓��E�{���Av�f�C�E�n����fq�2�\-g�_���d�L>�L�(�dUA�5�F�BX/p�X��	TH�#��=9!��.Z^S��;F���"�������c��i�M��ՓWX�!?aw�%�Nt�G�����Ҧ�������s�k(�ܢ��"���m"u�%��w���9ؠ�͏���]��d������	{<�U����y��20ţ�k<�A�(�dAi#:&�C�V]�@K,�ƠO��g����%Q��n��p^������O�?16dzn��8�L">p~�0��U�Ķ�ȃ��q��1"\yohǂ��+�-�4���pޒoϔK�O�������I\m��s?C?�e�#�i���M��'�OQ糼�(��v2��̲"׉)�8�{�l�0�U��ĜY���r�O#ǛwK��%�+�q���&�a�w6.E��I\����w)ݟO�*i��U�zTFO�0ڟP�nbt�AD8����&+��<[Ү댙���"��U��C�3Di�gVP�j������gF���/�
��z�	�����}�`�_��DCk>��3(^��4��z�#.�'$ZFr�Q�hr�����w�i��*����90+�H���n�=%��e��~�ro�k���k+� [��uy�����u�7qL�f@��1�ص�lM�+��I�>��}s��$�6e.���ś�@Ѭ�}���0��Ƭ���T{�V�ɯ_Qħ�U�ag�_u�/�G�B���j~�
�ZI*Y�lTQ��%\'3�aԃ;�)@����� ��#���%��Я���탴�x
ꅎ�(�q�l�$�l��u�q�'�g	W��t��wR+R��չ;�^��摫Fn,��TCCk�U4_(Qu�R�ܞ�+reD�DI���u$�jVF<C�DM�E�_�ʚ��dn���:���n�X�/K�
F�|�~eKRV�t\yӅ��!Zs�&��I�7նM	k����˦� z*}a�/y�#
q�K�S���ȕ��
F���)���w�w�R<����3�ޛ�Sx�Og�%��4�%��9�~�I���*U�y���ݪ�x.8��~�h�G?4,��� �o��������J���y踀�>W�����NX�t��=滃��ɖ�.�RnV~���7�f,?�JXK% ��}uH:�uv�K��Ph�� ��B�3L��Z�;F� ��D-Ѽj����n8|'$�Tg �uY��z������O��9��ß��u��2���� �w;i����u:;T~l��enw�Bq(T��!=WzD	<��ьr���9���9�/�y�/gA�#�����X��0���t`Ĭ��������軀����)�pDr��P5c��m,o�v�du�'�����B&ix�_�����hHL.�%���m�|W� 0S��ո#�1^o�%���jÂi|�$��u�
8����B޼7kagSN�`�
B�������OO�g���P�[ ^����BL@�:WU7��t�	��K.�{����W ��:i&ofrO�4�Ï�\sM�bez�� ��ɷ
��A�5f�<A�]�9��F\{�Mkv����R��߻���
�Ћ�����kO��$@�ڶ��M�K:�O$�-YԢ�7�+���󁏦���m�%̺��x^��5svibY�y�g���|�� <"4e�b6_Y�
�3�	:hX,Mi>���=�(͜��mz}��4�8D�A8���v�W��^�܌&W��"d�ALw�o��pQ�̜�ʩ�l<�r+���\�H���kj�ݹ1�Z�����u���;x}G���0���!6"hӬ��T�;ԟ��-�
�C�o����i�����]Q�m`V���SQ��<4�������O��1")����H���N(�EL����QJ#1Ko��]c�� ����hѶd�,���-z��J�3&����ҏ�-x^9K\h�	��m�#0 +�|E�sI_�}dA���3�PVpغ\�J�B�lU ��%���X����ln�!y�y��۹��aIU)wL��C���blik	��-��1o�9 Ÿ�)�q�Z��)�F�]�Tx��bld��?��8����bZ
�@�:��0c2�����^�d�}�#�6�Ew��x�.;�1�_����5��(��"���}sL�`�V!�nv��=NLL�',c�w_.U�6�C"tv����ު
K���"����&��f��:ʂ��ћ�B)��X�<8����}�{"uB��K����"J_�8���s�{�<�P&�K$��o��I�͓���2�L�Bl����87?;kPMo������&��)��3�8V���rE`��d�^!�H4�}鋝�w�v`�U?���ڠ�Ld��o�pݹ�Sr����S6�Zz���M�f�q�Q!"!A�r�.v�c�6\~֝����%�0�_Ճ2KJ�o��1q�G�(m~�s',�8lY���|�"��ND�h� )XtK����5�=��Z���e��������VS+�]���ȸ��X��;���Ma��c���#���2Pg`��;�ѳ�A%P�GJ�ͩC�hj��ٕ���vp�-]z��VC��6s6l`��%�0
�`f���E�"}�ɣ\�����Z;�f�ת���b4��<�Psʷ�lŸ����g��Fd��#�G`�T���N|.BN�:Hi���d(U06�J���dd����|�"���T���*�%y����ah�5�NdJ��r��0ͱ�N����-j2j?�R�SW�?�<�B:����f�fh<a�+�' �(�Rc|�7���?�/�t�M���$���<>\.,��b9~�C�d����]3*��d�Ff;��q�S�Y�G����i��tL08e����Qr���|��{���]^�����۽&��罙��K`��+wv�"��	,��#P�|j����=��]ǟ&fM#��<n����d"�����J���u{��R�M�\6�Р�<l��Qk��b��"V�<�	k�{iV!��5�D>����Eq:t���~��|��P~��g�*W�fgQ'"����]"�J�2ڊD����/��0qq'����U�x�)�I9�։��, ����e��г�� ��ǎZ��C�������$�05�a���[�\ȫ�qЕp ���`��$�ch'|�lg���K�[�Rîa_2�:�_}�)�հ�o��	�x=���K��y��ȿ���U��YC*V'�RZD��y���,��5tF�+-l�n���I�N~�'�d��S��ٜ>U��w�=1A��{�9�b���!��n�ֳ�?��2q�㫸�;�M�����a$�+���!�5���X����q6�6ZU�x���	3u���z���;@����hHϜx�(1�k������x��iPY�G-����M#��{6#+�+Y���	�d�ЌĆ,78��sk'wjS�/?н/GcAk[���W�H}��RWt�9�lK��H�nr�;;��=�s��v��'�v�� ID�p5�����I������o-ݿ`{a�!ȗ��d[�cRuQ��G^�ͬŗFςw�P���ݻ�0*�:~�T��M�A���5'�?�L �[طǨ0��(���y%ƨ~N}��_����?�#�u��GӨ�� Ix۷�Ք��O�e���BQ�0�VXYPt�=�-���_������FTܱ%ScY������ �Xg����/����E�ʰ�V9�4EX�?O�ڙR�%��	��T���i���-�ڔAq����U���mFV{y���'x/aW�Q7�l�xB�%��w������'���$%o�p1��6dK�M���}F#�?�:l[�
�^XY��3�WBm/p<_p�"�	6�>����g�+�3��)!�yĠ���
Ju�r�����{�9��jP�*4fԃ� ���&�@��:mp,̫��x�=1��	YF����_u��1ʡ�g�p~�C�Ƶ�EHm)�m��,e� F��tOMLWD�ȋ�p[^�B&��.qԀ�s�F�<��}����g��'7M��SE���[�6��U�����T�jq)�{qJ�7R�5|��)t��ꇗ�+n��!�<���$��TZ���O�t��	8��+��K�k���5��
����z�@�=<(B�d*ż�ѧ���r��4��jQ��g���^%�(l�6�-�8������E����HRD�����>�؈^ �!�� �Ӟ��R$l�t�V�����W��_8������c�N�̭�j:��ǘ8�lM��ʎ���n��0¦]=����Nw��Ӄ>]�t �G承���1�#���C���R�Si�ˠ�?�񞦆
�qN�c@V��zٍT��Fo.i�D�/�M�473p� �9�d�!�
*���������ݤ�1-������e�k��V"ھ"	�1�=���ɿ�#��B (ѹ�����X��;�$&/�����\�idVn��
Ygկ:� >���4wH�
k��9�tk'Ĝ3"����L��eE ����Pq;`�qip�}p�
M���\� lYO��b,����l�c�#��.��J�вC��k�A�KZ���!��v�OJ��5��g0#�q).���`��Z�����r�B�:}�
�Ĉ��Z<]�%?��J�&<U��A����mm��H�%��5�vqMqG��Ð�}���r�'�83{|2����F�k/&|���"�%����� jG���ٖy�j�5(Ն!�P���I��)����;�Yԧk��?W�K�-�������������꼸TJ�c����$�
a���HI����y��s�(o��|/��UTD�y7X�٧t�;\Y�v-�|D���"v��Od�v�^�o9�+8�&&��Y�����!r)k0�����I$����)�|ۧwe�!xH�$HA�����OSvYgwy�ѻT��^��5|ںC�oa1�[8�%b��ne�1��c����7�3�F�:���D�����'d���*�m� �ďJd��GtӮi�_��u��a�]�:�f=�>FSƑ��x)1b
9Xg8D�В��;��|t��E�������rV�2�����N��Z�|������zE�����1ɣ�9 �!9���v�/Δ�ӎȑ�*��p5��̮m�HX�q�2�]���[4�񗈖����������K�W�����{Ͳ��Ԥ��#�D#4���|K�Nz��KC]����U B��9a�$oJ���J�nR�}��׫�U���<���q���qYG!h$���K��ͭ���Ҵ9uXb"j��	�3�x���#Z��}��~�&t�mC�����`����:�[W��	�GegV;R�c&W.��+���I�,Dԏ�
�';������R�se���5��턴�H�@�\�����Sw����/�.�˴`�%����O��CW���E�eܗ��Z%)b�.�X��K�N���y����o�C�
M^根��NHJƥFj����1]��}d>�Byh@�%�/%�������A#���ܬ���G�L���Ǆ�E�J�d�P� Txz�����696�3<�΅frt7�C���ڗ����=i�6���fYꟴ�]����:,R5Uڐf	2Ъ�?=;]'���nA�6!5����}�|�w�s�<ɚ�D�:�]*\C6���2�B�@O
^]����3�+6�x�b����T�["�E%X�=�E��:}j-}?hPeI͸Q�@�+�Qzc���[��.�wt��\���6�O��#�s�"��)\��v2����!"Tk�$XN;��KoƏ�}y���!N�Wu]��F䇩�90E�HSzӯDB����
��bx���1�sy]�p7wG�lh:L\XFt��cG��0%0�· �bu<��P����]7Y'DҤ�w�C�(�_Y�M���x��rw���g�����$;���[9q�1�VU�lNБ`Y��`�@���*.l#�PÅ��K��r������螁?��^���Vuj�/_��:�HBlj�p$_"Yi� ��Z먔��ݬ� �q��A��X̶�@˚�*my� -�CW��-a^G���v���Zjw;�x�D�4�Ȅl�̸�o��籇�����M��V���{�#���s���3���̼�-9��NGs�G!��u��;�Ӳ%�ΒZ�m�L[66�Ջ0A�OT�����)E�WȖ6�/D#Ql��b46�{�!0���ۦ�	� ��ә#�[�S>���W��C4�!�BV"��߶�1ʈ���Iȣ��ZØ�9�������� j?��/�=���R�pMwOo���.Ż��A��3$5��8U"些����I垅-��6���PX���1ꉦx��Eo��$Q :2k��W����L�E/,�(?��a�C��d�jm��1��A26�fy��)���V�uw����`-��N`X$D��H����*�*`8�2����8ǘ=��hP�P��Q�-�cR$��мt
>�k��X�Oj4���
L��e��P6-���[J�{n
S"�/b����Dg#��z��M4.h�Pu��?��ے��lE��M5������Kʄ_�����L���
>�����0��N�~�,z���49��$u���#xE�������v3SK���3H�%Av� ��m�������ة�p�Ʈ�C����|!����i0Zw�J��M�y�'�yV�򽖌X��������,o�w=�Gе�� �	X%�YC�C����㈇�S���I�5۳�K��q����Eӄ������h/V	��B���6�m0f��3E2%q;v���Y��St��,Q���j='�͍��bO��:�"+u�|vHzꁪ2~��V"�G���~�P�Us����c�OF����X��G���)w�V�	1*�W&2�%44q\\"~��������@y�ȝ&�E�J��?�F��il�&�9G��sG�%�{�4(?����ӽ�4U[ۼ�!�gW6ﱨ��<͠_O�Gk�9&�ʺD�ʰb�g�Fk�:�R�kWq���=���]6:��3��~�?�Q��̇���y��ڳ�HX���^?)��"V����%A6R7x��9$�>��r���7r���/�XLX2�|���>��~�����<v �ڱ���Lٵ��tL�Dx7*)�	�P����y���M6y�P�1<9�^�|-%;�|\~�'P�G����?��͎�Ő���'��#�>SB�a��M��s1?,]G���?J��*��wafL�p���M@���J��E�&B� ��U  U>I��Gna��Py.��Ή��3�z?���{�@)������*��%����zyMV�m��O�8pȲ�e�LXE���p�m�(�v���qe`��;�'��Ϫ�K�&X,$k,8�B�ߞ��#.%�N�ʸ��	fr-��:�,��R�&_i������ ��κ��wP��c��7�ǵ�*�-�)��Đ��B�Ft�ƾ���ap8|����-�W�z��ԭT�h�;=�<����®��m*��q߮/۱>W���K����v�U
a0)#�|����P"�>uz��&����!��=U��r�;GX^�ѣ�Wt�I��I�J�]5�1�YM�@�h_s�F@�bF!O1����E���"��)DGP��A#�W���SS��ۀ���j�v�V�B�	�˯Н��Sz'����-h
����9���������R)~%V�6�����t٥ɉ��5���FBe�����{\޼g����b*�w���e�?����Q�#��u�%�F���2�vvy����Use�<	��	3��-�[J_���#�˂h:S��2���K��#�PBU�Z��ͻ��Xձ1���˩�,$��&mǟQ#>���Ŧ�mR�q4q.D
��h�荎�?�*$�6`2e_�ARoH!������p����G&�+���ꆣC��'t��=�+EΦ�x�.2�jpX����^�"�c��`�'o*�Fr0��v*!���շ�8{�i�Q�>��*]/G��	g�����B9��#3�M,%������G�=xjz��#����W�N��6x��d�a����W<�A9��4 �.��ڻ��e��&];�=��''����<nm�kۛ��
�yV��E:i�C��Q	XW[�������'����&T�a��,���s��_Y]�m��h䠶�7Y��<����>�ܘ�{�B��y������5?#�$+�#l������L�RĜr�3���˖=iq��`(f=h���#ޒ�}��A�0 ����s�y� �$�v�����(�πV�wY��U�,��GН�1 !�I�)y��kk�NMU�ĩ����Om!��<R��iLG|V,t�JF�״�ȍ�(����w��e��(�>{ 	�QU�z�4��yJ,��02dNR(J�S�,b:�n��cP������4�Q�G�ԇ���qhK�U�$���!��ٞ�R$7��gT��U���/���]"�/汳�EV��K���(+��S�Xv�!z�݁�RA��5P�IGu0zL��Ѓ��9,3cQZ�>޿ޠ6ա�P��Ք2�޲��n��W��VC(�ׯ��A!�[�i +����֫V{�)�7[����m�j�@.(�%ˇ+ק�7�U\E��O��&46��-�$�	�wEi1�x��9����y�}g�* ���������sS�07-�e�DJ�uz �Ͼ��_I�e&8�a\�s�o��hX{���`�I��'���ܴ~�գSB�+e7ʃt3�|(,}��f��c |7����������(�%֝A'"�l����U���FJa���T@J�[���k���c���z�8p�n��j`f��r+U~*�@�Q鰇Q�ە-����F�'wT{<��cR�J�!][>~ �����[�[���۟u@�^������H}����O�������Z��|h����r�} s�<�>χIt�gro��<u�����k=�%�$�L���b�;��AI�����B����g��X2^�S���"�*�f�IZ�j�ϖgW/N�<�B��1� G�>q�5[��6�9-��Zl���q��M)%4	'��r�
j���8w�!pCyZKu�-j�ј�h5|���o�� �:�ۓnp�}����%wC�������ԬnN.�2���(m�W�z� �H�E&�=��&�eIՊ���$�M�FŽe�~XY��T�d�6���>�T��X$������^t�[%KZʸ\�K�.%�X����VPyz8���0>M
*$��*
�*�j�����d2�#�-������$d�t	�P��b�&�5k�82yI���g;����{ V���p4�Ha�7�)�o+�^'�}��z��q0|h�l��Af��Oc�1�_"�Ysŀ-�,�=nɉ��V�Q�o���<WRi#�l�u}�0�XC��-c�l�u�c��b&y����a�ړ6tϘ�
7<�k��m��R��8no���c�쿘-��!����Q�����	)؃u����-����
����9��ˮ]�b.�\���bu�|Q���,.(3�n��v��r�K8�g��?��Z��	�\�K7�X�h�t�Ⱦ�b,�$$JA�ӽ�)�a�Ȃ�@a�
�1�2/9'�����2+Z�y[����`ĩ��y��p/�S�K����	oB���/ϵ�ءV ;�1�y��:6"�g��SBًy'��鎨ƖyXѳU���T�f�'p2p�u�Ro5
m^���P�bO���Jڒ�tɆI��Ծ}�G������^L��δ�I,�j�&��Q�?@B��&	��W��a_ߐF!�)T1�|S�� ��ð��ųX��%]�#�xU)aOD���&~�1�� -���z;��	1����K��מ����hf��VJ�5���U��0o8�^V����if��_g	�y��e�=�9��������X��4�d�����a�D�v:4�A��ϥ�O�����6��h}2�����i�hU�e��8��$ܵ�G"`܄������˩	m��������_���B�o!���E�^f���KD���_����q�\���P�Ƃ�/�1�d����~̳��y/�{�#掽3C!1�_z����)�a���.��d�u����́2}r�3i�6���3��Z��\���2`|����ARX��Iylkn�2>1�2���1�F�'�aW>�R�0�s�������|��:��NJj�&�{���B�[h:�����A���!Įaw�l�������]�?��K �J�c���"�B�����å���)�3K��,�a�ϓ%����A����s�p]�>s`Uԋk���ǈT�Ӭr���|p�Lo�Uf321����1Q�%�֫tc���f�^.�+��3L������R�+���-R�AZ�����w�kz����(/ps\��Ef�A���b�]xa'��Di/��_���"ׄ�3�g�H������|u�sO�+{m�}32k�|M��Z�@��9��8X��:d�e�`�d�i%��akE�;*�"��L8}��x/?�;��͟��2<��mq~4���jFF�T����7�YC�_Z����/j��ly
{{�����y,ҏ������[�x��fU{E��J[p$a-�MvT��!d*�P��yE�ezP��?kH6_�W���^��4BKZ	�"M��`�*畍�Wǒ�Ȉ+��yU =Z�<�Pɝ�r%��5Sx���[��V[��O�pO[i�4]�t�[�I%z!���0�<�n?��R'v���C�c�`�BTi�N����Ѽh'g����W�C\^{*�K���9��O�köFB���ka2���l6`�����y� ���T����.I26��f@Á'�}$-��	�E��f���'B��v&�ty�.��RK��Dl~F��h�3����)���
��E�x���$!�+���mM��zݲ�����.�IEifb��?�Rt�����������:��I�}.eO�
�C�u|���g#�J�sHzzX
�%����x�?�ǡ��q\v=����B�f���VP?�
m�b8��F�4f�M��(�5�戳�H>�"7��MN�g�&þ�C�����!�!�LI�7�|�$�QOD�?�Ǯ����2ٞ�>��O\�-{�<7~�]2t�깺"�j���`�`�1��&�>�gB?sQƈ���B���C��&G�_^:`	��p?h��� wdzlU��}�|���1�W���h�Qt��H�qd�?$f�K�j���<�����G�y�,ߞ�,��[W���`y�-!�G!cS3�f�qˢ�|E����9{V���*��Od9�ތ<(|]I�h���'�Suj��ɲ�����~X�"��ƙ�"4�ց�"�n����7�����Ӕq
���$Ī���܂�����
M���
;ܬ�L�UU뀋��  ���$$�c-?��M�w\�[:�y+�(,q�
�4���iu���=.2�m�B�do �{����o���'�N�ȲMBޅ�D�g�����6� t˒ @��-�҉���#�L�p���0�q�����B��.l�1
>�Ŵ'��@��#U񐍕F��6~�w����
���=NRW���pI� ��ޭ���<ε�7��(�~��K�:t�Y�ɚ/iY���w.?�O���D`�"<�"�W_�$[�x ��)z��<�:e\�s�Yv}���>��ؒԣ��(i!4���nȟ����¢�.��r�%sSσ[�u�k1����oRgL�zs��&ˢ��x�~E�	�]�eN�u,lc`ip�M�6��e�QS��$�N+M%�g $�%/�����:`��-ed�q�`ŌM�R����_�5�̲R�^2ӏo��òi��C�u�}2�=N����� �i���4�Se�-�Y�B| ��K�:4��� he�S[�	̚���
������^}��q)�9<��k��vYF�)r�Vp9���7LUݡڐ���`sKk�7mVV7��V���4]��Q��@ZD%���-Mt캯Lg�%z�l����?=�����M�g�=���ƿ=S~��e�j)�k�]���o�˨䴜�L�����fy��� ��_��3�
]�؞�M����i�@ ��PuK���$�5�VK8f���>l�8c�hvTyOF?._K_$x�����U �_�^��X)�oI{����_�˷>{3��\ֺ���d�o��1���#���G9��0��[P�Ʋî��I��HN�R�[�v�Ө�	�>;[h��]H(q= vk�<X�i�K�AµU�;�9�Q�2v�0u����wX�s��?�Gq�?�<jW�:8�n?�Q8�;=��KC�$�l����گ������ɳ�����5 �k;؆�C��W�s�!9d)_&Ҽ�>�8�|�G|TD�	�u���IA� ����Ž��&���p��Gh�v��7������Jg��h�39�'^���A�!����ĕm��>8`��6���1�4��Oy�-2�S��L,�9h��q� �$j��l��$����W�����-�x���Yb��{�:��b�� Z!���D(�(��P<U��EB�g��>B�0	���?-�M�
�[Q<�_�o�Z{.C�4je��!&�mk1��m����ؑ;��;�¼�??x_��b&{�;%���qu�˔a�IE�����>�o�1s�.�.�};�L=�������PQ��ފR�w���x���������ķ�l�/ �ch@0n����/�����Э`�ׯ|&��t�e��'k�)[�7���D�hQ���[��a}�&���b-��C���9�w�ș׹�8���{���d�!!��N���ih̋
�F=9��O���*��~3��aQ�� >4`KL�x�`z��+`md���V'¯�Dl��OU%���f$�G�:��
�)�A�|h6(�>0x��Z��וwF�0w�<�Z�3�Z�]�(H�R��Xv�)%�NӐ���y4�?B_[՘zVY�Ze�0q}���W���"cu5���r��gJ3û�7��]ot���3r�0de.���\GXD�:N��$uR��� �(��)�Σ
n]/I}����f�����1gw����?FM3Bw�=�N���9n������x����G�8�SM��;���0����0M�Է�P�}�=�J�C���K��C�+3��j�߀�W�l�i*��򹷧O_�ȇ�Q��wi]p6�Ո�`lE��6�m�_�$�G�i��D�k���r�����H�5�B? ����.f�5;Q$k����ь�d��������З�5�䏺\f"���!�`�k�h�'ko�SCI���Mp�xqO%J Q����M���jIo9@Z�`��^aU�A~�{�mA�?'��^���1�v�g��"G� ÏOf���HP�o+�q��r+JJ�%UwWrIo��m���a�J�i�ۙ���Q�`��]���&Y��ROy+	.�*»�ߠ�M�k�����BlV�UqN`��8�w";��d���.V��=;]t{���H��+U�@��������|�h�~$�������ٖ`�s��yw���	��n�$C1"B{���F,7T�Գ&����\N�s�{�S )G��O�p���ի�S�#P�I0�Pxa$��.�,X���,�&�E��N��v�\a�t�&�~=���!i9�V�1�q"�L���-tb���е=!�˓��D��� ��wF&V<_�KC�(J^4���}���[��*�4o�эVm�wd|h+d?��k�Z�jt�?f��m�>����b���2sK)-j��k�N��@n�C����E���S2R~pV ��c
����Q~P�k�W��`�g���D��&�č��L�b��!m��`����1Vp#�����3�� �3,�n�|�Y3)w�
�+FwH�lg2�H��eț|����<1^�A����Q��G���*@���dա��m>)8ם^eT��Й�C\����/C���Y��5΢!4��r����_��at�.�б��mE����Pz�<`o�Oe�قǮ���8���ء��X��V�W��<T�ĭR�����0d����;`
���?��ܔ���BHƕOr72�*6Rz�6mx�HD��|�~�����_!?%zN�ǹ����u�2�(����x	ٽu��Q/����S�?��ԯ�3B�
{��|Ѱ����)��H��+�
�tmii"����´��H�ݜ	��N�0-����٭�R�MZ���F���c/X�#U���d�������q�.\�W����QƎ�9�
�7i*��TY���wxP\��S���7�V��9 ����þ�A�yW��ݦy�H�D_>\����T�iD|_����P����i�D.Gx�vR(�X��/�I?�����Q�8r0n��m(�:֡��L�jZ�'���w�����hP��b������:9yd1k�T��M�� WM��E��/+��=(��N#�+�!�کm	����<�\��p�GzΰD�F\�m�x�@�L��[�h�4߈O��;	Z=�����N$����a�OX��JWJb8��5���CxJ��c��I�����h��h��!6�������N�s���L_t�v%�\R2�}D\��
��/h��z«�|�.X�Mp�<[z?��q�;��	mA�o��u� ������.��p�ƚM'�S5PX�ŚR��iDVA����C �"<9��jc, ĩC��ld�qR-��$}=��m�z��V8%Y��w�aX�%�+�.a�غ��V�Ԩ�«o�O"Qll�O��I�f�_���O�'�Ӫ��Tʊ�i����%�iB�^�"_���سGg{e�	l���#m��1����t0=�8�&3g���˽<�����L��ע�xOs���!�%=F\j�W��SUB�N8_���fS��#��ʌ3�b3�}$����H��]z�=����~T$��%���i}�0��GN��g�;��>���x��8\r��qWԥ[w)��>�z� �K_#���g2H6v�����L�g@��u���$s2�M�T�M<;6@z�uF��⢮���D�'V�nK�}'&�l���Ct���/J����9B�9��̤��� �V�H �B9�{z�-�Q�p{
3��E&��1���ּdw�w�#�5#�^)��7�̫��;�D����m�h� �8��ۈK8�ABp��`�4ڮ��Ub�������!������۠x���~��%a����濁�=4���6�~{���V1N�p��k�t��)�,e�{0�Ј^�� �4�Ҫ.!���[�0�9B�OtP\h��ji
�Y��jf��C�5�tia�g�6?`�Aq@G�A���r2@>m�����$��p��A0n��rh�4�0�1�~�����i_lPĂL_�6a��4ΩC���ɟ��R�R��eO��lt����f��V�ߞ\hZ�7m~W�R�ꦧ����'\�~�p�-ѩ�^2o��w�J!��:aj'��/�2��c"Z�_pҩ�0͙bl�B�+��Mjw�b, 5�!����J�!�h r>��]��O���&Ҳ��.�~����*��p(��%����ش ��Y�
"B ���=�`4��#VD#�������Ԟ;��N};��f泝�a���b�F)��I�뛻ʕ_h���i�ͦ���χ~��e��?≺^,#{���|���*��HA���7@l}Jt��� �?c�]GԉH
�oqe�H��T��o3��X�7
����I�����p%����u������ԩe��Ya��7��V�7*x� ���)�%3%ů�>5�3� �r����G�sV[)�Dʬ�P?6�N�x<Xe�UI�=��ȴ�ʮ-�M����X����f�+ғCXt�q��$F?�����e)����ֿT�<���=�Dj?��\d��6�{��SHD�Һ�e`�6�L�y ����Z�:��4�W���	��������w ͛��s��5J`���I|�ף�K���E���QO�H�/_�	�D}�Ƒ��6֊jEv�e�������d'5V_��p��,��%D�\���>ZH����F#�r�a��^	١4��k���!�b]���#јj�r'l�L!�T�K�����ҥ��屫sT��*� 5����+�Bv� ~hFe(�ː�ｲ�h��Q&�C��7vd��?>�!H�����Fkw+��/��'UF>�i�-� 8A��xW���ԅ*"�X�.�>�5�~���"3E��[8]����΢p�!�-�!��`<�Iͯ�zuը5�1�AG���m�z��4My�f#��oU�y�B�"Z������u���.���� �8��:8 �Vic�=���c毘�k퐰�X�*Hkc���b���0$A�X K��n�ـ��>���t�Rl�1�R���}M��m��T֭�~�����4<�lid^��:`���{=�Ko7�}_S`��E��7.�;�d뫌 � �Ɓ��XݱL������v*��^P�~$�Ui��F�S��v��,������r��W\M\S���a꼹2�L���s�l>]1Nr��͈�E���6��|M+ko��w�W݆��R
+_���e��@e��o��v8�$f&/c9LBG�k�n?�zKP�n0w�㭥���5r�g�z�\|}�5+js���$��o����L�֊��D�;E�-!i����;~� 3�<Q��/=9C�����~�d���`�P���^4!u�i����+����Rw�*(�U�,E��Q�[)[)hKb��\p-�d7�n�#��3�/k���s��'�0��.Oa�D�an���o�c��i�Ž���L�	��$��3&��ƞ���t�.�ͦ�)�U'�Z�1Xgp�(X��l9��-�T�Ø��S�\}o�8�D�d�
��Z�m�.�pL^�NÕ��9��*I*߰-sI�.�bi����Q�30ԲT6&��B�j�=��y�� �BYM$ؑdB^�0��l�!�Ule��4��o��7i?�pe��F;���_� w{З
Ian9�7ʽ�~��q<|MrXih���^���q�+"�a<�'eيn���Y�%���@[� �Q��sUp�@O	���BuB��^�D�k4����8+zķ��9z���%f�Ӱc�Du�L��`3���@m
7J�FLes4�����$9��n��p�S�x<(��4h���i%Qg�3��Pšl��3��K �ŒJ��o���#���p��:��w��rz4Ih|��5�ۺz��^�I��u��-��R/5L�WP|�3�*x�JH`��������'AA]�p���&�X�di�T���mZ���o��I�(�X�Q�)s������7)s5�?#����f�)q�A}�4��t2i��t��?��˺���H�#�Z�ߏ�϶A?<`������)�1S�p����=|\�ʞHZ���� �ZC�⧖��-��4����d[k'�#�}ii�� {�"� �#џ�x�NS��J�>��^��g<�G|=�)A�E懢㴜ڊ��Е�zB�u�2"�VH$�7�/V}1/$v���"Ns+>x��?�Z�.�ʚ��J���lu��;���?�8������V�ʹ��;h��W�7{�4x��|ynl����������);�sg� H<�GT$	d��<f��1���2������H�a����U3�v�(M�=����Z�*���j��)�׺tZ���� t����<���Ȇ�v@��گb<z��v��M V^t�G|#:�;�v?�3>���Ԥ���dl)j|gܞz�o<&�]��]�UWu��N�b��Z��ƌ�_,�32�*l��3w�[v��`+q0F��D}�KRC�H�l�,s��~�����������5�H���@�탷�#d���ߖ�M�O@���X.�k%N��L��N?��@@OH��8$�z��߄�H�}�=V-��x�P��ם'�9�.GF��cV�m[���S��<���[�n �".��m�m�����������M�z�"1�}ʜ'�>��X�Ԓ*DgEL+qD�NL�ߑ-s�p6����<�ѻJ������GL
1@T�*{[��Y�������]t��5yW0�>�h38�i]BN%�pid�_�U�����T���6h%��^񢈲�-
����Zҗ)zD���}�QLq��-�o�2���QOaz_��Cq��wf"�Ҩ�Ȕ]���@e�m_	V�A�!ڻ�#���.��^[�7;��&�F�uyv+P8���g������P�&-��?[�N�9��ׯ����>RsƎx�dԥG�?ơz��/k2ߦ��no��? �-R�01�V���^L9t.���=S�FUt�<��"#��$=�5�(J�	���KlΠ�� ��Ym��f���fY�7����7�&;�a�b�y�B1jٿ57��<���P�4�T\�G��U	�b��o�����!�ؖ���D���ωu��M�D�r"�IPtQ��ac4�S���;o��L{:|@$1AJ'�B�`}�X�	�vH�R��LEL�'�� �X��9��o4/�,�A&Y���=h���_�7��Ҋ�9��ݜ|�s�������Kz|�O2< ��Z�L�b�],z�9�^��<T��i�z���-kIgq?���h���  �D���+ด�;�|���9	��gE^z��P��|���i^�'O���]=a�gz��Y�H�^/�y���4���W���z۸N��Z��$	�w ��,̻/���;��o
�3dN����t�j����:�m�<�k��D���E5���������N�$�k����kz{�S���U�m��#��V^��|���a5���(:��%Umvn �i�@�xʝ����K�zϷl��� W֗�z%1`����t��;g1���ku�ypD��k�u!c}��0W��KOݻ��q��z� Fun�OBq6��)���|Cà�B��(
�_آ�1�RU�iM�i��Ej{I�G��;��^i~d�_��פD�Q��^���I�����!�:B5`>D�m����||� c�_�:]�t��ڌF�?F�����ʂ�X��Be�=�8���)IУ��uokW�~�KStY߹��E�����xM;�V��Wʿ�����V��h�.H����y?�ާg�DȚ+_�QXr����(�!�1��#|t{�7�T���.��'?M�7��W�˗���N��nyKv��П�V� 2A��֓P6(�9�f�߷�C�V��n�J^.�^fz!��3-���*_Z����>V���*�AtM;n�b���$�;�޴ъ��S�-ߐ!�#}�@#{|�Р���y�1�j�Y�*��%�p2w��1���dvڧ��bM	����j�f7%'V�ܦ��b�x�m@���e�K��������?��pW<�W��bF�J��50��^���D\�"i��&�sM096;�nf��z��rȠ:�p�!�s^X۞F�.�$���L�ͅ�5-I��8�1W8�D���Z�Iਘ�Dn���?��~y��;6~ϟOP�#���V#oT�aY���U�x�Q[���wY���]�XF�.��ږ���)���  }��3�}g�����<"U)�,ӹrh3mݣ���O��e�<PQZf���z��F(љ 0@�V��]�=�>��Oe$s���,)5��y!�?�ķS6C�W������i7�@�`)ǘ�K�<J��U��(�REx�4�~��� .%J���2�/:��c$�˪���s2�k�������g�����/<8Ӽ��l�m�+��}��o��ԤUop�q@�oF�R��#!�zH�v�S��T�u�N�d�Ruh�2<̍ ���&T6u��&�e����
�X�qӟotQ��k�$V�� |�V�sp��=C��-�-�4��9[�D�j
�֏�<ʆ�)�j[[�VWEO.�ٵ��d� �X���C����n�xЃ��ف���xu�GR_j���Zݳ�mV�'�mX4R�ր����oD�o}о���|ra1��s#�amrq��.):�Ddi��u��M=A>��T�cV��U�iNj06/��A�Qޠ�P�B�򛰆v<����,B�p��]7�iL\˼%5���Q_�`%8?U� o�۷�#�	5-�j!��j\2�F+���Q��I���?I�L�UU8��Y����̀^�=��\��D�[3c˗M�����@�R^��Ỷ�Q��p:��h���𒦧t��yVcx~�0q������j�@u]0Z^�`y��ꩂ�5�ݕ�-㠕��Pn�����e���>�/�|�+�%V�m���O$�U�tr���z���qZaŎ!B�̂��
���x���Lfma�s��?���bU�.�W�����q�r��r ���&���U,|�gڲ$��G2������D\��O��6����mu���������>��k㒘������m7����|�����7 ^/D�P�hc<5�*�Ȗz�jy�G�K�%��z�u�a �:�dG�J�Z!��q�v�b+���ֶZI4}���'�B��w�F�E���R�����G�P�c�J��HI���=B��H��{1�+�Lpr�>/Թ�I�p)͹���>� ��
�e�w��@cs��_&�i�����|<��1{@�!��"E���8��V���b��^�pyF
3��'���G��{�L�pO�"�
��C�mF����?:���c-sh�X�����*����襽�����������ӛ��)&��ZC�H4$��i�aq~44 ͱ�v���=���`;}yX�.r2�[1���+欬�?ʆ�4�׵��b��g-���m7b�0n�w�vc�RͿY9�܅�Q#Wc��	�a)�����S�{����������@y���P�z�޻լ�9�WE"�*W��*b!���$����Ya�aB���K�,X���ǖz�n� �V��@�1,�?l���)������i�c<�'T� 6^�[�h�Q�6�f��X	+	£�A�5���ӂ�/}J7)⥷Q�ߛ`�\V �_���'�v����Ju_�m��3�����#>{��+a�':Y��iO�LK�-)5�fP&��wT]=Jx�4l�L��q�n���^�6��`�����f�E�{�4}��Z~�q{�3��J��-QCc��{�u�I�ѡ#��
l�J���Oo]�Y�/�K�J��*�i��`m&g(�!�S�#��)c㝭C*`"�@�l�����2;�>����:��5[�5�_����u���hƙ9V�]�))7���]�;lf�~Y��HbL$Kg�Y��Z��}���5��f�ME��_5��?V>�U��B�1Qu8��d�^V���&�3����ڋ���IF.j�t��b�޾I]fX��űH#d\Ϡ�c�.w�=�YT������l�Ia<�$"x�h� �a3�~-@��Ҽd�<~��j��>w8���0���B�뽖.6ق�Ǌ7T��Q�$5l���k������?�c�mm ����K�uz��w��_�I�ǓHG�?��B��cmF�L�9P��g1��dz��%�����է�� ��Db\|l�����@~ ^�nEh��+��`H���`��2o�� ���B$C�n���c�d�����
6s�S=a��#i�I�� ���[qL)��l?Ŵgr�ϕ2������uԦB��GK�����	.��>�6���e��'}���]D0R���\Ғ�s9i&�}0�9#�ڵb�jREŃ������ϐ��T�E��\y,��+�Ud�ݟ������
χ}v�N -�?����*��:K�h$����H�_S `�B9�R���5�9g	}OJ��A�}V~������0PPd���7�K�T��yh�l��DuJz�C�l��@c� �>w4Zl�i�q/��R9/�qÖo���k���>+�d%K�g�
F�n<���p��n�:8�����=cߓ9�[
.}v�V=�r�9]��\U
�������$,�Ε�t��dBC�*�)$�c�{;����2�܌>�̙���ɑB��U:&�V�C��z�|�G���=����hH0��'��dԾ���a�:��vE�S! �j�'j6�ҝ�8'�����B�ܸӅ-��=�y g�QL�س*��E��x��,x���/ 
���Y�#���Ӑ�񄇬"���D�H�<����9��x��"ʇI�he!)y�pd�?7�d�>�26�#~�Τ�����J�E�Iއ���զu?�!�3O�UZ���������!�>�hr^��scv�����)�"���e�vR.F`OW����j,Y��Y�y�������d��OQ���[���Q�w�u<�OX��:�3Wj@���&/��:DD\z4q*�,P������6�%��_n�R�{Ƽ�~�>wO�,3,p�VǍ��"�#k����}������[�1�y���D�#�hyƅWH�"b�
����B�2����c��5s�8��/0�� �Z�A )���/��R����I:|�^�{�p�{�gV�25����@���LR���c�ܨ��m5�p+��+q�ˊ�[��l�W�r&�����_6z$�7I�|9�fa�����oX|XKs�9��
�G44 ��+�|��>C7-]!X�� f�N˂| �[v���Gc)��b�ݹ�Џ)1M�i���= �T����a?��j��%�+5��r�Ȱ����*�@�/�������t�����_#d SI��j��|�����<F�LXc
w�5_6�j��'�'�RKD��;���)��gt��8��-�J��t��+\���	/&����)�o#�l�����ަ�HI(j:"���hk%׸pBF*��!�۝��7��܏��^8o.�&2�tp���Y޺��ʛ "�. !uR?eEk�$�3�U(+/Q#󦖽��_�B6���S(���u��LؾA��[<��X3�C;(֩vC#��T�F�W�)F�A�A:���%6 �{�D���4<���w�S�V�(������E�6c�(���C�H�)�ɏo�X�HB#�5��X=d�C�Ԥ��+s���	���#���I�y�/X�%�,�s� �F#|/D��3��U\���������_�|�_�x������.
������-�YM�c|̿����/z�.�2c2�>	��p�I>�����d�/9, ��Fw;}J[���8*�^��SJ�YR�C@�lj�3���~��E_y����0�,Mz�:i�I�!͝V�L"�o�8A�K��	A��x�;��I�@{�'�gH�/���-oi��J�r?-u~�b�y�7�9��!�6�K���mM�%�<�M�  ��\���Sr�s�<�{>@�A���*�Ʊ �v�KG-h��J��0u�-�ᇼ���1��N�-�e�5oO���
7�����p#���96�\��}��,��Aq��}��C�DT=����Ky�.�a�[�w�y���V8�bfto ߣ��/k�@�W�Uqz����� 7 @�$q}��ޛ���^`���4�3|�:-�mw\����j���ggN����n\J=&x���/@�;�S��oY��laσ��%�x�����S�!� o|)EH҅��A[���E5���z5*�S����
\.c�')l}Ѧ�G� ����.�ᅣ�\����B�X��t�:˘>������)�K�*n謰j!��8=��B��j�ŸDљ�5魈���LR���T�pky}�m8-hrt^w��Y��%ru�����*��Kmʶ��?3�+�^���?	�h=����!E�d���]ӭ���wS�jB�r�y�G�d�Pg�c|�8��p[%�p&�9��l�謶�9t:��ĠN|�?�D-G�_����d���EE*��Qn��B�"�����|[D��[uY�8�D��]�`CL�2~*|VO~�<be�:K�Kԁcg�z��]u�qųa�G,:M�y!��@ī�'�Q�gM�Vl�AVL(�8;���Q�Ô�u'*�~ )�$���osd5U�9��$ء�4��v���Xr�k�Ҩ�����[	��� �����b���,���p��W�s.CK�_�2�V��e`Y}WG����\2��J���d*�݌e�W=���>�{b�4�Qs�Z���X�f746 x��[B�ێp�ȿ�@�A	8�h}�NMh�����t%���n�;����\� O��mɎ�T�b5�V��k�HS�ۣ�/݋�e8��W�ļ2��,����YpEԄK
�6T��j���d�{4ζ;��k����{*A;��|-=D'M���Gλ��kL���Β'���3�g��r�T"&�Rq���3��Z�����"z�}ȑ���A���Zu�]�<ߤD8:���I�E0����❧�W�"s�p��+���E��j�`��5ٝ�T.��"wOyIg˗#����#!K\7��fjσ���$�O@M|=eғ�Kn��.�e�iZW�jn)~U��e�I����Z�iJ�8[�t�h'G`���=yX$���5��Ϗ.��<K#%�D"\s�6�m������̟��>U�%gF����?�	�z���;�PW`���5:��8�V�	ٽ��(f��RF_�,���j����tx�!'�|��T��G�4��Y�i�
��
�(��#3������ᾮ��VΤM�\������	��%��'��;��z�l��.�f��l� c�JY:~)�x�;��.a��ZǤC%�_ԃ]��D<*�Χy�§�>���M�����$�R���ֽ�֕�$�s����_+�š*��H$ce�Cnܻ��&���|h���Q��s��h��e�rԕ�����=���P�&��ϕ>�'��S�r�9���S��4y򘉑 ;i?VIw��E��j/YIҧ�  �w
�yꮲ��1G�F�������5[.=���Ľ1�ث^�%7�-C>�Nɦ�d�N������#r9Z� �f
S�jZ!]�`*��cz�
U��arӮ�*�#�,�U�	9)G:�bcQV¶3	4f1�Q����o:�R��OM�S|�g�֔�
]'fԏ6��e��m2 7i��Q��C�V�����sS0Z�.c;hf�ů'7Փ�tON���lS�r��x�v�!�MM� ��,��ǌ��,�p[��$��{��!�thM���x��ɓ�MR
,����vS��}�k{���L%E��l�w;xT{��;��YH�)�D����g��K�ټ�aߜoi��n��1^��TK��ym�`h�^��̘�]�9	Ι Ʈjk����=��T�� i|PR_g�jc�� -#�� ��`���1�����s���8������"���!���X�?i��9��E4�V&ĕ��j�F��ƭI+p�2�@����jL}�-oG&q'|]t6�\O�l��p����O��!����D�wj��J�si�p������UB��YI]������tS)O�!?�*���	ʙZ���SPn��-^�85��1+ݗ9�A�.�����cO�+�
&{ݧŪ���oH�{�]�,�Ki�^̣�7�`�����R~�3��Q���)��Y�q�����m�rw]O��ЛwHё�\�!���:`H�����b��;g�������Fm�~���q�q!	g��,\�,���w,�p1 ��cuAe${۾��#in�L%�N�k�~NN�l}��k2�sZ=���{˕�!�-�����V\�z����*�U2�L�qj�v�0�U6ބ7Y����c�mc��V��
��e�I�Q� 491g�;�R��y͊�� ,j�e��û�źL�D�{K�����GR�Q˴��M��T/6�cy���� �Z�I����)W2r��-�p�(�]�~�����(2	J8����5��=��kʻWk�6Q��у��d� m�OIo�,u���q��Y;�U;���A������f��L�Wiz ���`m�y�Y`�.f��`�G�c�'��!�Ԑ~e� X��Q�)b'd8wz<1�����6��yAb�p��ߐ��ѽ��*��C�'Mq3�1�J|7��jН���k�K�A�e��v�=�(2�����fq}E4qF�w1�0w+c%�г�͝��ȅ��DZb�,\�ZVR �������Nt�ǡ�_�t��4����
�ӫ�4e�$�6��y���Ğ��O��@�Y�D�h�\��������%ģRϫ�LB��T�1aW��̨*��@��9G�F�m��hQ!�""iU�-60&�Пf�~<�>ފk'd:1�U�=S&v�2Դ3�t�M""��ޛC�{���x�7�C��E��P��Y\M �W��{b)��}�� �ю�κ4���5�_Y�^�~�4�H?j�O�.[���Ob��{f*�f��(8o��22}!�Fn%=�C�$����	/�W[��}���
覾�3w�;�]�_[ڰ�[���/��`�R7��D�����
��{��Br�\ݶ�V*bh�Ѳ�.3!��_Ҝ�֤������.�Z��.�,�y[�x����x��i����#�r�cr��%��tL�1�+�_)���}�uj�kI@���y'3��t��������w%�R�]=�2kl�8<��m|�� �>w�,oN�����	It.8!a�)]��#�ᄗw��Z����[ذ @�I�N�9�hȨ���V�e�Yx[�8驼�z�u�!�.��� fΙ �b�dh52h�Q���Ay���yW�]��}�}ց��儀g�&Zh�.���������֔��^��W}��'�ITk��$�)�KSQ�=�s1���k�L��[@�����U\1^��r��pw ̸����M�A�@���~��2���=�r�bn{C�A)����6�
~�	������Cv��M�����C��׎I��]ثKJ��je�_bi�a��<Y?S=W�-[v.���/c���4�6���Q�Cui	�Py�+\W?}tu7�QGF=ҏruԵ��M�����C��|_��ӄ�/��|�>��W���`�y:iw_2c�����^gwu��\��VH�U����?[�FS�����?��4����R	�%*�y���nR8�t��|A����;�{�5�uZ�A�o����\�Y�&3+m��,�kj�cd��(8�`d�����3Q��6���$p�f�v�C�������n��^�I��!I���I�tg��!"!V�B7=��uH{�_�ty	�Bϒ���7P�NyJ��D�_� D�{��F��ƕ
*N�����b��=G,� �gU%���P#.���r��_��3����p�L���b��.7��1_<MO��ܷZ|����~�;i�1��liqcK<31��ݐ�|��ZEْ4ߑ@gAQW��P)(=H�{ټ���@��e�Х�����gP'�x�'����3k���Q�sb��6>[k'�2�7�����#f�v�ž9 f�n|��UǻvU����ݢ^2�m*�qOL#洳�p>����l_�׳�s��H�K+ztA5�����I1'ｽ�1l1��h��L���(F�R@ۿt�I��h=����?s}��.������Jo��*X���������]�F���뱑�������:S�B��J�x��~�bL�c�fP���_��VG�	-��>>^xN�n]]���0�	�M�|�Q\O�ˁ9L�mRδ����h�vK0��7a�M�m׏G�/��eyh@v��ıp������L' �T$��T�L���5F��D���W>4pS���Q��~�����b>��-hv��c]d$a�
��Ƈl��kԁzG�<�.b��Y�*;��k�H.��g�2,�tX�(ƶ�����N���\����X?r���C#���� �R+k h�'<]�Bڛ7�/�Kw]���h;.^{�},����bqj������'���H	!��K>��P��;^GȔ�@�ď�����o�ɥ;fo�Q�oU�j�Jq�*�2�<�Y���b#S�w�|,�������ؤ��\?[C��M8�%��4�{g��������*���b�f�=SU�J�VGR���\ӡ�� Ѕ�[�i�~U�2�$���؏�of~�¯���+Z��j�����A�w^����������J��ZpE���\���e�~fl�=p��vêx�K(�C#%砃V**���ט60�d�f�w�ؓ�oUi�*�`28�H�g��D��t�d�$�f�� �mD��]@b�	�a��������y:�+����O�c����Ȗޕ�\�@��ª;`+��V-��U�|�W��c�����=�6>d�ϗ�v�0��<���1�5MtV�rT)z�ǟN����& �F|\&����	T�v���Py�^�թ$��`U�[�e�s��7XӛX��%�N�Œ��
>3��%:�}X}��x%w�g�SP�`bC��"M�z��}���I�'�pI��� �(45	)>8�����)G�Q��pb����'$ܮP�T�x��w��]�R'�]@3_V�����%����'92d@=pq�e^a^sr����v���}��ڝ�~����Z?k܎ȁG�џ3|E���}s�͹ �+��)�J�J���RP�q����^2��)y2�����fHH^)Ԗ�5�.	�Lt?�������H�9	U��8�9�������8��6�p���M��֋Z�X#T'�����7BZ�&P��^�4h2�( �ՙ�2H�eK�~���6Cr=�ӓ*����xE�#���s�,_~rDv��T
�}-�S�"0WY�%�0��=p?{(:�Mha�#�DH��T&�ԮX����&A}&5�r��*��}�l�	�8�,�ϑ�ܺ��V5���}����X`���^��ހq\:s��L����Ќm-�'���a�W�"�@��Xj�0�; 2��)d�^�퐂�u��ZI�a60��i��±�	�qo��?z�F���cX�w����t�oty�+��c������^�!�~�I:I��O�E�D�녯�dբ�ވ�8��Zh3.5J ɀ��腕��H����H�%k5*�K���6Wh�Kb���� kP,�' ���|A��*�3+����6�l#��Qθ
P�:�\)=�M��CS�����řW�d�J�_��x���xi������{��'���<q�-�2A�w���� u�o��K�a` �i��W> Q�*$��i���G�7ς�1c'��U�3�g�j���/JGuiy���?������g���Hm�7z���G�,ʑuO5�2p;kQ�;�6����b�vb��Bd́����EPr� >[z�fX[9Yl����փ��]�p􁸉�#�^(cd Iz�I2�s�:gQ�����a\x�z�-z�]��I(�t<>���ʏ�Y� n�)ΩPSwc[��SP�ά�W�'S�3eVg�����מ��AU	n�]$�_C�'<tGܬF���� �Bq?�����84'f��hy���D��s�7q���2t^��b'Dɼ��a�����-��M� ���N[�Nz|�qZWy����Z ��	�n�X�����<�,����7熓�X�;��0��Nh�$��EW����S�;��3e`�v�T�TU:��||�;&�-�!�i�����$�M^J�`���5{M��������w�d���)�Uu�g��m�����Xox�-.6�/3�]&�GtQ��$�N�
�.&�J���+Ĺ�0F��<)6�J��s�a�f�$�Ȟ�E}��-�M&�ܭ1`��ݚ;����M��X�=@G,�k{��VA�@�+��H�>�b=ݩz��z�Y'{��|���t8o�qM5�r �%)}�l�ќ)�)8�L&aN*����<���E�"�}��  D���oI�y��H����Y
=��w��&��n�bCiƮ�pox�D�_,��b�I�UnmM>��O�+H�⪺k�������ĐO0��T,��/���S	�4OW�~�Pi�wt�.����E��z��+P��u��䘦�x��àHy�q��[�" �^��w�5\�[���J�h�ȞqN�`��2.:���q����>�����R@�C��|[n�B��z�:�潒��8p���<9�d&jE7��	x�0��2̪�(֖i��Η�N����M~WP������b���)����:���D����㳵4+a�W\�C�%"$���Z�'e���)d�"����>���g�ћ��6�[t�)�������hK��.VW�+rw=u��}�dD���@,��yd����V��t����\.���t	4&ޢO�s$���kg:��)(�M��S�y�H���cO�PaԱ����dsrP�&��U� 5�����G��?���h�F��PY�u�� ��Ve֨|2bHq%�s�1Hj�}�|j�R�� 2�Lc~d��)|tަ�`�(�|>�G�y�B�Nc��>��#��۸�E��֩����]��� S@�2������r+� k�%;o�,Uד�Q	A������XW�D�?9�x�[r�l���b#AA��ùm�R�P���з[3[�#"䠶o��f�S,(�`-�����2�|�.�����0�yh�>�V�
(F�n�C	ɱ�<:�gVf��[�e[J��侅
�Yxr��/�4���ϷL��EM�C�&��k9���Ԥ�ǋ�h��n�����G\Gs.f-x�{�ܽ�2�5,Y8��MGF�"����|��t��}����k<��go`ǧ9� 3gs�D2�-S���6OLy�F�q��_z�6KӝK�D�A���4�� @���)�Z������0�PD��u��ڬg�z�xu�[P�������ُ��,M^H�]5놟���Q��-QԋYZ����D�&b�T��MP��mۑ��b�a�r��s� ���.���Aa��f����	wj�G�U���c�^=JNՑ�|\UQ�N�D�'h��-��J����-xh �FX�Ç�A��[���\*��O4��HA�@Ĉ��H�}�u�OL�;�3W2�ADPA�>�d��H���<y^�:x�H�
�|�B싉�Z�%m[I��x���M����*��sV�cu^	pkӲ	Lx�����8����Ө4c���

B�YEȗ�m�H�~��q��2�)L�p�T�)�ʁ�S�g��������I�e��VǾR�%u4�����E�1������T�4�:8�=��u����l>���2ʨ�����zE,ĸ��#�
�I���C�Τ닧�M�n�|��X,� �Z�3�PU/�1��?�ǖ��'Q�� ��>o���T�U�6��>Y*� ���@"��Pyy�C�F�o"��)G���	�'�8��K�CC�\o�Xb�Le�_`%E��-Pgnv�*��Mm�\���x�զ'Po�pB-fpR'�P�\�866@:��p���f��g�=m=p����<����T�"���S��b��V�!Ϳ2��q�����_ ��^h�o�b�m���Ȉ�T�S�bF�B�)���=.$'�٠��i��*�����AYֹ� 	�������;�H��W&���lc�����1-��J��Ѽ�����w�+��	S	�}p��\��ZC|\��
���Kc4,�N2=�*��KAYa�����0(�����eвs'��NM�����$al�(>M	��xbTr��UE��j�.��/o饂T��E�Q8��%��Z�%�Qf��'d�
>��D�7Q�v ��]<mU�&�\�^��/n� ��t,X�A�S�x������]6M���4�)o6u�^��H5�J��ǰ�����f�3�FԦ1�C��KCj�3�V��G���+��TtYE�r�������
�|��+˾2)�y�Bh�*>������H�iن�����O`���X�.�B���.�~>$��2�d�&L�7�?��D��
�X�4P[�����������`�{%\Р��>�,�G�Bʡ�*`W-��.����4��*�4�@��_2t~�'�ohEs��������[�ZT$��i�D�6v��_��n 呁��zo��(��N3ǜ�Ԛ{�t%&���W���=���p�])�jɠ��^VP���\ރ2�d%64�\��N��_^q�j6���syƸɠ?7�y�"A��h����f�Zo�'�܊	�Q`�\z��YtI� q��P̺b	 ����`�����2�O�td�qcS��E��g갔�����T�+�M.��ob9 �� ��Z�u7!O.�ך$��h��([��ͦj=IK�B��%}�pU�����V�RK8�fw�����0�w����4T&�4k�	��f����uH�Qn�Ʉ��=+�� 6~��|����Hv7�g���d.]H�K��dZo�����1{�Wfn���=E|�k4��\�;�}j��i�cd�d
v��� tb����^r9�P5�[��ځ���fA�U'�����	=�J���qe�J�ԡ��S���Z�mt^�u��z��"R��G,��;R�ꛎ�G�I���5+y*=Z��W��Ng�~���{�"��Q�[B�X:���OQ0-�꒥��&�����F�z����ߌ���`K�� ��̐mG��d���<3�� cj�T�gj�ŜՊ�a�D�/���_���aڪIc7��#X)L��
����Vs�!��� �׫�rK/Cp��/�f�v�V��!QG�d��Ry�����8��,ځl~��Ʃ,�䁰�s\J��q���_�hH�_�mϙ�O[O��t��d>�(g�=���%9�j�2:�Ǳb�F���N�ՂFU��ګXH�(�np�#J#N+wٓȑ毙�����π��[X�l��"+)�4�9�ZI��Æ��Π�D���������~���.(��p�QZ�GP����Tˈ��L���n����N:����Zrf�F�B����X����".w�n�G.ы	(^�č���l^�|BqQ?�_{Cit�[�\���8L�֞P��~m<�6C�(ŽT����!Ȟ㗍�C�	Rt�p�R�g�43�w��zJ�2hs1+������[��3@l���!9����f�Z�v'+:D4.����NO)�[Y��xv��������+$[`\�T����dy=�z�eѭg7�R�ҳ*�p��0�d�(A�
}Cl�XA�ӟ��%;%lH� W�� �5eBٷ\m��Qh|��m�+���@R�̴���o�p� ;͟2a��4/ܛ��ϴ.[5p��y3�m�Mn���z����ip���������h^!��_�yVR�n�tG6�8R�_� ���+C��@Ylu�cإ�YUՔ�B�]x[G��|��@���_�j��~�*�����ĥ�p��x)W��sdUc�~�ri@*��� ]96�t|:��	=��a�v�}�)��p�h��ys �4+'}�0�e�(�zw���1O��j7���I�;b�ya��݌�6��x�P�d�ٰ���xV�����&���{	��(A��[�<�$yj��u!����Iy'��!w,��F��_̃�n87)�h�����>&����K.ǎ_���Ѩ���AmH�5�e��tV-�oZ�	Kܒ���i�/�<-�'3NE��a��>q4>��e���Ä���S�gtX�Np�|f(�n3�6����a2.9���[&�5�^BBm��o�Qi�	C#�$3�8�9��s�R+�b���p�o�!jK;_��ƻ�ug,�^��ۅ :�H�)665����2*8�%���Mq���j!#9��/cQK!��M�K.���K�� ��	U�?��Q�Y�8-
Tx۳gq�|���z�"ԏ�'�a�%<�ᔛ'�=kgWs�k����"��7��*�J�&�ی'2��xC��j����"�c�d�HQ6,ӏ�鉘�-��^�q��0.�)�}��l��_<��rNS!A-��fv��D��cQy'1Ol�-+c�J�=g�L�3j��P�?~�VHm(ڙ���ȝ�r�Qxt����{	+/V��U����~�HB�0�и̾���[�#��@�,���]
��B*yo�'��"�`L8��5J�{=�	[J�H����9�cokx��h�����P_D��4�X0I%����hom;�x6k5U�OQ٥C�4rڅ��a�+�:�ç&�k�i��N�3��caˈȴ���c�$��l8��(%�+�^�@/�s�3��ڝ�pk	����ڹJ���td��	0;��e�k.kx�rvDG>�x$v��+��utxjwvr��/W�p�_�����Dt���V��Wh�lH�g�x�Ԕ�h�-�(��VFϒ�j�����h7�r��B�ف{���C����X�>6=�u����Ծ�Fʱ�ț[��������X�09ȯ	���������n 5�`��F�/����ہ��1�n�Q���sX[}��H���v<�sQ�&$B<wD��0�`ɩ��v�#��Gsd�BWNMMX$�2|&��h����$�ij ��w6���^��#��c=�|��՛i._�r��k$>Lv*aD�o�]Gq/�!�֓�d(_�G~I66��t�q�^N��!�K��.���CT�ϝ��8G-����:%���A�E�J��1�p�l���J��� ��@��f��V{D�C��>$�mY<Tt��D���.M��r�K� >4���y�X�Nkcva�gf�K!�6;h�'r��]h���?�e�i��K��}�hR�O�a��гW��&���05��9�ՙ�,�z�M=(V��� |z|�i�E��g-M�R���Aj�K�o�z��Ƀ?Z�(�`�LL�?	)������3H�#�������(X��V�.!���[�L��O!�$��l�h�d�#��V��	�����
FT��8r	hE�|z�`����	��y�3�D�c�g\�0�(]�FS�
��y�0 dF\2(����Ѹ�}�V=�B���cGv�8��D~�����2��-�K��VTo|��QG�C�3G��qN[?�Rm��zҶV@�K��s��왿�8���?��ټmmq,[Q�+3T��#�ޛ1���~���4��gQ��u�=���A�Dd�У�3^�n�:>&"��y�g:����KA�YqK�hC0�XҰX'����H�*^�:U
i���K©�)�n	�­�Øy�2�B�RU��J��T$ɜ��	3IRp�5��C_�CX��B
�UO`��I�볝:󛳎?$���Վ-m#��<8g �[����RL�f4���p�Xq���>&<���հ��=����닛l��֠�5�u˾7iWV�P�e$r+��4X�!��fpe[ܞ���Ԫ��57l)��_pK�1J�t��c��'<c���P`9�tJvZ�×rY`L{72OXd��p��;��ֆ}U6�]�-��A�E�Kҝ����?�z�	���]O<� TR���Y+n<�sRu�'�Y��3m��c"�w�o�۪��ޯ�$�����`iA�6�­Jl%��@d�6�9U_�Sg���48���
�}�>2�=���es�3��9�߂?M����,6�H���öQ�].Y��ܶ�,�k���(ʅU.A%�-�����	�\k�E��v@oZ��>�����.BJ�����]��F��W�J+\����0)�P��6e�ns�0yjy|���ޯV��B�un�H'�I�"a��8�u����Twe�}Y^rL�qu
hx�����u�)�[��#b�.N=�]Nc�N�f���d� 0.��	z�is3�Μ)�Ї]�"�5 �[��B��߁�2��%	խ=C�����'�f��x~&�^>���:��]BqwF=���"c��n`/0�ct?~.2#��(XB?��&�{ʈ��P9��\���q�ɽ��-�㺞B�kw�̑o�R��	@��^ 黺�fxդY������,}Ѓ�����!�v2-�|�*YM��l��Ϥ�l�]Hw��B/�E�����/X3�d&g�&���z~�J�~�b�f�u9�#�TP����~^X�K9�ȅefb��sBg�9)���ѳ��sC���,�-VR�񂽘N<J*@k�-�$�P�[m��_C _9����drP;���ffO�����V�6�F������
�dj��|��[�c���`�ļ��,��Sw2s42�pi3JRL��a��)m=4��ֳ�2Yv��j�R��WC��܋]^\<q��+���Y�_[�b�w�MBD~�->��ܚ�Ɏ�D��1~@�J��`�Tm\�Xurj�������l#��)�֪�&*�-�(<�#-����`y�46��/`W�T�U�~��.�;C:w֠o�B�ʓ݋�A���戥��?�n����56M�Y�Iѧ<����lH�o���	+É|4�3�ѬP�Y5��SL?b9���>54
3�ϖ
�13�Z�鵙��v�nFk&.��oSح��3��U"�2�+m\�`�I乜�������ї�����l��u<2T��rg�$ �q��y>� �%�ܴ\�e�߃+���
|���'�/ܞ�Q�5'�9�������E���Vۗ4��Fe�a<J4���p]w��@Cr�9�R���@8�e����('�p�����d����l��a}�E�x׽�ΆF�^٢I�o��jy�o(��I�T���`!n�7M�wlC�w�9��nq�<`c�mp��P�.�4
l	yh��&����'H`ɂ~��}7�r�)�W ����0����|$/{`r�~�1�t4�(��*G��)JJ�0�ԍ�<��?�pv|+8��F~�ڝHNHk������RgN^�E�;���u`��`p;��+��F}E�V�f��@��lS�T1<
8��K��bf}j�k: (7C�g�V����F��}@�5�N�_$���E����;��16�ܸ�w�s�;�y�HY����Y�)F�nKk�{�D|�S4HNZ�)�Y��)R'�<������uL�M�"[�A��L� �b�
�ySC9�<�ʄ�~Җ����oI�H���,T�)���Q��#�S�,���2������h-D�ѻ[�OA��fX����3TM,Et���}�YMH�W΄M��5 ��a��^
p?�D���%�	j�2�x%ν�*�w��`��86N6.�9Wx�ފ� �KH�u��5��]c��&����I��|��@?x�-;����=�� P*O�@ZKxEnߏ<��R��9�Q7j&��@I2�w��Z/G��̈7:�5��(�ʊ����h����]E8>�ܲ�}��6vrBsf�w�X���+k-|E?��r����ڛ`o�}a#��B�!1}s^��4U6����y���%Fr�1R�\��SO`Q��)��|Nn�/���my�dOҪ�5ħ3�X:����x�^��e'=Wd;�Ct0�d�j��䓲��Ig�ap��6�i�p&�KO
#�}�g"�#J�`�4?�B�~�A�O0�Ơ�+��n2Z_"����O%S��0��sB��/��m��Z$�W)&��1"ʧ��h�r]&��.��·����{C�;��C��P�"�ZA(K<�o@&���C��,��E��싑2�\1���|T+��������|<�1^[���� �Y�@�*bv>�3��� Kz9$����̻ ܨH�6N߃)���=�'k��W�幮�P�K��~��W�l��*�_?M<��~�Y��%g$��0���QU#ʖޡ���[7�>餟��W|���a������3w�@Zϫ�0���̘��9��ڥ�zK��:�ˬ�*�
u�[�՟9n�u�#d��� "���?һ�����J[�
�H`�>ۣM>�^����]4�W77ƀ�W��T�*�z��� |�@E�B]�+�y���!���|�J`���EO#�}V�k(��J���C�U������0�P$f}��]������P�~0�x]����ȫ�0cy�G�*o����L�w �+R@ @]t�G��F�"R���'v�� �J��t N�u��:E׾�,��cT�EPZ����E��82(����ߓ���	��҅%ɼ�ӱ�w|MS!l�lXo�m�f=�(~���O$kB-q���^A'T�M��rb�5���zhv���Q��s�E��4��1�l)ٗ��P&���F���Tx!����B�O��sN�n6�ڊ[3� $H��s�e�BQH/�57��H�!9�l��~C���&~Y�RF������qo1f	p���f�`g�s������U��j���Z}��S�eꋭ-�#���A�_�6�q|��hL	w'WCۂo&� ���BO��@83;���i�I�*u�z[K`�񛩡o52
8�vU�W|�C�`i1��Qy �?���r۫�,�7��R���!�*R�@�����0�O������y�˳ltI����4B�@���}l��LjpIԘ�d�oRC�Q�p�*�E��("�M=��%����G7�$�V�u@|�����$�
d��W�`�=x���[��2��ȴ`�4�&4��ږ	ժ@�(@f�߰����J"���3q\��O߅4_w�ʽ ��A7���D(�C/}��Mi�J�b��uwsFP�u0&Y�GN8�1���T��Ȟ�P��H�"mGV
x���Gϳ��u_"������� 0~$/�i��m-�)���Ť  %%��{�'),(��@)?����	v"䫯H�,�*1���t�DB��{���ߴ�#�Y��E�m7�T�OfE�u.����'	�aĺFnMF߿�ߺ����o US����~��ǧ���:�]��3�?��c����7�?�����(Pw/��X��r=��|o$i�A�<Щ@X̳���$F�1ݽ�J�b�/��Y5�&��Ղ��3h�|�Qyan-D�T��G5������ Q��B
h���J���C�\�-�Q���'f�%�P��+�4zkS���M��#6BK��ƫ�{�⊡1�����n���Ps
�S,�ni�S�8�/'�О����xF�9��J�e&՝���n�QCN���6p&,�9��okF�'���
�̾h�SQ�,���p��K��c��W�&�����'Z�N�Gc�d�=�qA�P�B�����f���
܄Ig��)�J't�F5�s#	,�l�l��ָ��
��Z�W�D��3�FTQ�a.�0��D��`Z�ld�"*���3�ݴ�I6�?��w�׶e�9��� j�u@3�%UO��װ~��$�?�S=>�N
,�L�_f�FY:��?�y�X_j�NA5���Xu����N��-����+xQ�D�Ж�,���g�m�t����;��%�=�������|���Ъ�s�LM�ې�1K��-���!������Y� �J2�M�A���`=iywHX#�N}CZ���|9v�AR�-gBe�j��Q�ܛ��|���p��򘾖�!I}�������$tnS��'�A��~�i�2BGM`�$u�2�W��ƅ
�L�9q��9��Y���@2�+p�̙��4�T��h6LO��Rj���^�bT�;��U��Ì��FQ`��ƈ�xxזQf�-���œ���+�R%�����[^'��,ƪC#��Sʶ�9��:�Q������t �M՜8�W��n��_��
G�D͔�eׇ��0��.4�X���Z��y��mCL��^9S���	_�U�\j��-����\+Auƒl�a�A,
��J�(�l��pQ��]t[�2^6X|Ou�J-LPWE������-F�iM�}Z��#P��.�0��b�X]���{��~� o߁��g17��CA&��m�S�δ�[Ѭ��r��?����~��t�9Ѧ �V�.��T���an�jK���ɹe��f	�O(�^:��R�7ޚR���{E]F$A��զ�JGy`.Y��Ll˨�f�№�V͖��^6��Կ���~�� ���`(/Q.��������C}@5�;��r/DzDۙ���Q|�[u��y�W���!F2��vG���1F!n��Ԋ��sCޕ+ڏ%��.���,Y��#S������q�f PB�x� ]�ě�{����+�Rs�ˏgMɀ6Pl���Ϫ�R=P���t��^+5�*��y�B����-� |��J&�B�b N�H����������l&~D��B�P�=#w���%�b�@�:"x-�-�|����P�h$�0=��;��<;PøzfV�Wqh* [��pwA|�4�nI��K|�`�D9R��G_�о6DS�K^�v�"���	�_�R�4_���adp}�4�I8<dj@UNy��U��l�����O⧷�A���6ٳUGj�I�R
��g�,Ï����Z9a�B����z ��kY�����0����BQ5)�25�wӖb�͆uU<��Ɠ*	��n$WǓ�@���pT��5q����t�^���`bW�xח��a�������X�/���
�9��s�_�7��:Z��^ݱ����\x����L�?�f�0�J~Ł]s�{a���X���:��?w��T�B(MoL�U~�~Z+j�"��|� {-1E�K��Lbp]� �/�A��׳)��o�mgǠ�������%����qC��A��*�N`d4�4���tI��k�/���q�oE%$"�A��F�ʔهfw�<�Q�fU
��7T0���AVo��;���<�e�K�M�L��c��I'����~��z������<��N��4�3�R� S7@��T-�O�=�k�[��|N3�������QN���y�����M��m{2"7����r;�~78��[��x.���~ZL���S��եp�(�j��[Jf�
G'� ��ǒ�3�c�z �d��L	Edn!��bޓ@�)+�MR��.I|/b�������y�5�b��Ӥ��$��
y�17�k��h����7(x�f���n��xщilW��Fn��9|}��nS���U�Cn�d��i0hjSt�;�~��,q��'TN������L���aWnF���N�9�#JU�&�w� Gdz�����!K���AE}N��/��FC̦���+��͑�C�Ŏ2�	��c�]�\R��~`�5��>QU����Co�`d�X̒ ���c
C"t�10�%��x�Ҝ�\Bz���(M��9�渤!����D>η�R};h���u���+$��He�ޡ���/�Z�"�UPN!3�(1�4� ���4 ��̑�r�h�3���ߟ �r?L��Q
�Ȕ�گ�۝6e���ҹ# �rG{jgq
1�_u�`�}Y�KT���>ڴ�']}b�`V�M�#��+^�B��W�P]v{�OK��y�����i�8�r������u��0��e��� .�DfN�ߌ�ăչx�#���³��P�Wu�WvthSS���!T�hX8���!��޵��@%Q��?p��-��A�xU�'��4tJZ���'0F��G�"�X! ��P:\t��tPM�B_ZHH�-��	����I��`VOsZ΢�%�9L�"�W�w�! n\��s��Re�,'[�p��v�X0�t�*K�YȠ�����X>��R��w2w+�v����[@�h��(�)=f��E�Nڝft7K����K�~Ƶc�ɤ��ZCƂ-��Ԍ��Q�b��H��'���	��'=�n�&�j�{>�M�ʞ�U���c�׺/A���p����Hl����EY��ϐˎ��
����_��l��ת� ��dc���j�q1l�:���~����4���n�Ed/KD��P�N�T��4������R����G4�Ik
����_œ~W�?
����w����� ��&�i>F�$���i�(`p?6%�d�m���/����"���^�][��'�z�����1	�>�����_�{�w��Qsn~@����z��7�j�}�%���|�L�|����#V~������{'T�q3�BҜ�aUi�k�Pj��6ntäJ������z�BG�!�%�FT�<������b�g�+U�L'��[�y���:��|�U)Oc��}�� �|��r��UHۙ��� 5عHU�{����N\A������=*�&��Q�����˓��B6��$�ٮ?=ڏOӳ&� �p��}a4�)��S�O$��F���w�BZ����#�})t��ܠ���ҙ(�_���m��sk	�	���B'/��yV+6�rP2���S�����s�p5~9L���iE�!j�5Θ71t<�b�qKS��������+@���U.�b����#��b�����dT�K��`eo[�)��o	e��뮤���Ga1$�cC�C��&�=��m�(>������:�*��:<6-)�S#<(Q;5���FE�C ec�9��D9�U����֓�+� �E	q�枂�{���e*R�8ܲ/���2I�A4j�a�
$��Xq!�����w#x�B��@�B�ω������,u��#���.*c-�H������[�!Eϐ�0�n#�PssL���O��ጯ:���-c���a�(��ؾcX�= ۈ>��T�o�7�F�/X��_�U�l!��'�g#R�JW.���3��u�)�7�\<�*�3K/�(���8�r���FGK=!�g��ps�R/}�F6���i���^<�&�!e\������s���BÉ��!��b}=� U�Ie�#��֕��#�����*�~{}+�S<n)P
Ϧ����qa��c1ۏ�@ڿU�N�?��°��!��.2*��y�zJ�k�W�Ĩ"4[!�f��f�BR� �rх������6(�KNT�M�}� �� ?3D�5���\��ޑ�$&3�����2nf�O�_Xp��c�4�n�Z�9��N^�F;WXwW�ڒ���46�6���1��r0���+���X=��p�}
U#Ķ�E�k��A� ^{�p��ɕ�a+�;��v��_Οޔ�n�%;V��`j�'S��a.m�w�7��C��y�<�w�--�)�ݛ\�{�4�Nm���Zv;�Eo%D9Zu�	�BG=ޮqn����i�E�������U��I����6��t�ʏ��6�K���<�x��j�9�p��Tښ�ǱK�\��
��,�L�L/u>,��$(��f��=�A'�*צ�Q�I7Y���ҳ�c$U��2�h/���J�y��n��2��NWM�<v8"��Vx� �/1�%�Mf�����a�N���13�J���yB�k%����G�Ԗ�Ò�x����ȳծ�Z�C&�������\���.��^]������g���ɌQ���L�����IЬ�$��R����� �X���Z�i!�w�j7H)��@�?��� ��b@�R��t��Qb�����-񇳀�B_K�΄�������dĶguTh��ڦm#�S4p�Ϧ�m�Z����	
�0d^�L�6����
������%
�����0��̒K�=�&2TG9�ԣ�� �F�����П7j;%h��r�c��2��ͩ��A�xo?E�6[b޴MƼ�ۼտ���p��B�Ю594ǭ�n�>`�e19�͈������JK���A�%9O/;�FNl���k��d��\,��?fq��w4صi��[s��7omF~=\�B�֏��X�-w��^!��cҫ���L�@g�f���Xw>f|�	�,��Jĭ�e����8�}�����5N���ۺ���±��H�M��(�6�9{��$��*��-5�����Y����h�8m�g��Vz_"���C?�y��<*����Ţp;~c��I��I%θ.<�W������=��Қ�N�����`��ykT��Y�<���z}#������0��˙�o�('9�
z.}�*�rR?;�
�a�D�uLB�Tu�S%�)A�觾�s)�Pp��Y���2|a�\yI���`܃LO�����HR̄��t�N���C���A��ɸ��ۢ �b��=�>�0��l������)OawIq$V�ϳ��pXJ¬P��o��<0}����n�թݦ�r�ދ俻<�L�/�욳VE)tR2H�d��s��ὩZT�����s��Rr��K�<�34^��#%
(Bo&^@�6��7A_Ε?X��c�4�����1"OU�u�����q��U��N��4������:��6��H�@�(��Иk܌N�������� ������̓�/�������c�r�Y�� 	H���b-[q�|�k>�N�%F����"d�����Q��M�к�g����K���)n&{o����=߀�4�+W�'��� 6�$���� `A�3�#h� �L�5g��)т|���R5�OJP�$C����(�Be�lyy��qoH�|I*�4��o�nƌ���F��3����P����d�%�y�o�~GI��Kj�=����UFC�a	 �7ئ��X{�P��{��ay� ���	���c���z���0�sj�dh�HZ~�ͥ��%�pr�{2	H{���-u�ʋ� kF�ݖ����p�L��v�h���p���
(�V�C��(�C�1>of*C�t4�+i �� ߏ3�V�9=���i��U�v9��u.���m�){H�y��C[?]����ijU&�f�i��t��X���7�����`�	V�]f6$m�9��NU��hP@L�R]����#��I#�(��8�u	|@�g�פZ��k`�d�%�=z�Է#*m�f9�C��R��Z�}ۅ�Bt����{���UZ���"m2zqUÒ�"!�BVK%\HY�1Hӛ	�l�yFd&����My�/���1V����77"k��+�*v�>��i5I�f��\r��At����ڒ����f���8�SB�B�:�$��w,�a,�'eV+��`7)R7� B�����2:����s3��sfܚ�����p���A�����>�� ��K�&l488tP�%��wqDG�Id���k�^g����:�rC8%���!�ޒa��|�z]���±�ܙ�A)�GP��9�W6�X�����4md�������x�Ei#�*�8�����lM������d��ŧG.3��ɡ���5�pĢ1T�h�z�/a�����:&�[�o>$CT�XH��NC�D��L}���[��u����ك2�X9�q��0���@3�΅\��z��R��嬨XN�H[�/�"+��S����~�!��ֽ}����5��N�c#"_���z�x<�M�X>�{�Lc����Vk��u�n?O��d)�˙�b��IA�:b�����`�2{�]�E>#�4����dAE���k�;,�M���c2�6��(N�ʶ]5�ӭ�þ�]6C�~\���0�T���c[)m ԉ�������QI#��4��6Ub����z�(nW�5`?^Fo�+�#�T���
=��7��Z���F��%x�@r)ɰz`�/w7�_���̴��jzY\1~��K6��?�six���9\��|��L����� ��6�����)�������j���<e1
g_�m�9����e'��v�����k �����U_��4�?���X�z��p�V��\h��Ҁc����<$f��~�.���78�[�4^-��N�1,W��	�O�<Ƭ�п(�.����ꗯ�f��v	%�k�ƴ��M0!{�r�z��ġM�
"�*��[��r���H�2�)��$b*���f>����ÓRP���[Mi���_đ�8��P���j�d�Nw���U�ud<9�G��Jϱf��D���3Jk]nO	w�r7�r���J���������ĺW��2n�9 i��@��n��ѥWdr��Q���j�iՋ���%v�����6,v\�8�����V����
�|��pԭE����_�R���悡��p�MT�r58 ��/�!��������$띋n��=AX�Y{��Olt.@J"T�Ik7��#Рu� ���=��Z�2��2�{:�9| j�N$�H??ZɞF���� 괯��h~����Sм���/�� �%w/\4��ޮ���(n��_�4:z7��}6����a�b�Ǐ���L>��U���X������
K�Yq�H���.�v����&�����r]T~Ò�p�xo�iw��Am��-��Y7Fɡ
��Y� "0��'��7*���7~��ú��:G��]u�)��� .X� o��ڏo������\+��^ᱳ��)��s�$����Xx��������ED7�$�՘��"2�X�B#�s�]B�w_i��ȧ��d�q X��T�~��@��5��豱c���xE_4��o�a�V�uƹ��(gX �T�o-���CLy�7��.<Y�a��>y'$ �bf^�.N!v�����zί^�7.�OL#��w�Cho��/ w�x���'K�0"���P'����cFX��^�;vR��-~�n�����M�����Q�āY�k9C�9�2J�E�CO�E}��i:�x����d��f������4o\/,Jw�����.QrAǈ�ѷ��n�r;�]��X5��F?P��e��g�82���*Y��2��=�Ubq/���~E�W\>)�N7���dȣ�+֙�~n���ֵ��f%al��#�zW�Q�=Jও�y/�E�_[�P�-��fÌ�:���ޓ�3!�֑��C1fLV�L�h&�e�B.�'3؅�F����n��Z��3K�O�H<�X�$X8�w��挗���ƣ����z[_�s
���ӞU��MH�,[�ߋP���n՟�8��{�T[����Rd�$Y	\�ӳ���A�|��+!��ĳ:�hqԽ�p�4�2?���L�h\bdk��������YNj*v�	r(V4�Y ��h�*���bV�Lp)y��H�yݬ���+��l�J�R�.�A���NdU��;_a�a�iiOУh�!�i�(�2��g�M1�f߷-��c�u��!�N3$���GT@�M|�(�ױ0����s��~mu��^�w}Z�@G� �y8�1s��c�b*D��zU�|�դ���2��E�A[	st/�}���|-����)F@}�ݭ�pt~�s�h�
�c����l�ύ@���pTV��9�z~���Q=��e�nh*��V�J�����l1!���$�Dh����$�J����P���/��-�9̵���R�����.m�����e��!�Qk(��=�Q�,iaI�K4�H�y]y��,�d��O
�}YDCc2�^�I��fWA}�ꀢΚ:@8��N"\/4X�v�A>[o���H5�����5��_����<+o~m��씈Dz4T����gh�.��+����^�������uL��#�)`n�3���y��:��� �p܆���	h�٢�Ui��V2q	����-���G�:�jPa΋9I��#Gm[D���a�tS����Y�4�U���A�>��=h��~�4o��u��s�s�Xѳp�`��@��l�ϑ�!Y��g���ke��&	��%�U�~F�+uM�O�s����>�Ge��l�k.1%6{�.��Ȧs{Aa@Ԗ�L��&Q��`z�����h�~F��"V���� ����3>����A\c�\��D��r#Pr��~jP d�>�l�4G�M&�T��ʌJ��2v>�*N���͉���a�Cnv-qJ^�9�#�na/�'`sq����#�S��`b���D�
l�oE�.������A�W-(I�9�9�s?���?9��681L��ѣG}&���ۉ"b���d����F̹�Y��"�������e̏;F��,�i����Ich:p8��X�[+Y�˭��p�X�!�Nw�;!\z�:� �ho�#^�
#�{i�=f�Q.�'���%W�n�%;F'Q�2M�1%��A��[��?�w�҈&a�N-m��N��¢F��+�������dʕ��;f֐�JD�/�k�=ZJU]ԀB���C��4�!��M��[ZŃ�av:,+�͌�;^c��~��n>������h�ĉN�[�l-���;,�pei�s�]d��g�xա���(׀��<�d0T����n��7A�B��EH��|qD����`9�=p���]���Z>�p�7�ccP������}��7�N6�G�Ԓ��/c9����<:=�?� s����sj�Y��P�ﰷ���R��� <�]�,�����oH�r�ã��Ϊ��c��%{o����b^	-=�Gg��q���q�t�@��/yl��9�7�D?&ջ�+Lm�c�zBH̓���E6���� ���i��<T��U4�4|*�P%B���x��Lp�3�:��Ž��K��X�Q��ϼ&��E��519[qC�����s���]r�X��s���Ye6�F�=��'_.Yf���g߷J�UA'@������e�|�8Q�[&�j�M�����p���e4�y��&���A�-���'	��G8�U�� HU�:��1��ҿ�j�r�N�9���3/�h���+��睏-���(�h����΍N����S�p��oc��#��5Q�XD kѿ k*6��k�9�h�;KÚ�m�m��N(h,=��n"���=�VH2sS>��H�]W�P'Ț�:>4�Q�e��0B����1�TKy���"��^>8F��.���^�*��2=D*�:���I~,j?G�&?��?���H��2z�Z��Q�(U������$Ļ�y�m���nd��p͛tqN[*�R��ZR�%�`}��mxRS�]�b�~ke�� �q��-��a>QB�>Y������>h��vy���fY�.Aj3��+΋�) ���e�G_��wKQ��U,_�ڃlJ2\j9%�
Q4k�u��@Eg{cJ�p?p�6��$*�Nt�k�a֞	=Vt�Vf	N��.ѫ-Ь������y+�{�ϣ�Ȁ���mk8���xW>ɑz8�� �)��2�>��o1}�=k�;g�������аY������o��j�j�_[���!�q�j�ii�]����4���x��X8��<޷�<�~r��Hؓ�~��F�6�� ���f˅ф�˝����N�5���2��j�B�Ǉ��D�.;�ݕ�1X}��m��(�s໺,��Y3� ��@j&6q8	�k�u���H�m���^)$��ԉ���J��+��%χݧ1�jl4��� "vv�Y��AR�DKX��4��%ӏ,��lM�)���jVw�O-!�+�	�Ϙ
q���cè��:迓6.d/)�.|��Ê�9��JMn>9z)gN{t�~����E��9{��z@�y�F&0�y��ᨎ3�Z,��M�P��v5�7.�t��O�ĥ����zE����9M��p�t��@�3�^���4������E�t���I�	���ڋ	���P��v��9o����� Lx :mL�8�Kk��k�+�$���$�q(����껁���S��A�y\ �;Ο��NV�T"�m�����"]5%o$y ��D������Y6�@�ׂo�a٫���e��jk�4;ǉ���_ϵ|4
g��O����@���,��XB3b�!��\���P�����6�u�	�L��X�5F��R�-A���$#ws�q�����=^J��l-�JG��m(^�k���8��b���x_A���F�J�Z�N9�b�[���Hv��q'U2��q�;�ATQ��
�	$J�t�l��m�����A����`!�"���5����U���r[�4S���Sj�'�S�5��]���wc�LMt�-��:�#���&�]�.5
[t�Qo�N�,��Z��` ���RT�H��aG����h��������n��������66��r��	z03��U�m= u������� �vX��7�!��P�t����O��pm��l�n���[�0䒪��R��傣��֫�+ς��)X���1��t�����^��0ryͿ�sp��<����u�az�	a��
�֊�������T�Ӫ��OƜ3�sʏ!������G��$k���V��/��FA~�Q�!aS�Nʘ��������C�`�s�8U��S���4�Tk�ĝ�?Z��9�b��}��/Z��x����!/�^�������$��j�0\&��m�/��G.�� �*�1�#e��8 (je��R�<������r������2`�ڱ]o��J��=�}������"K�|ԩ6���S>ɨy^p/N5���{Jxj�
�?h!F��#�����|}����ӏ$.t�qDG	�hK�gU�|@�@�$�	5�ɱ:s���G���9|�!!��[�GMf�{rP򴋨L���az������cg�6$�-�H���y?(j+��L��u�C��?�T)��m���o���e�%a�B�nu�t�N�c�pR�OxW�R�¸C��yyζ��!�����Hyǖ�+�n�ԙ �`� ����8�i��x/�<j�X֙�"+��E�Nv逹f�>w�ҩ>��[��?������o>+�	{(���A�P��Et��$�)모�����}ۑ������F��W�p��
����^��@J�
���+���PV�ीq������H�kh�5��b*�N�l凛������U��a�w-41���+�#�������X����� a�-��bVµ�<��蚒o�V�뤬M� �8��5���L�1������M�#�0�Mm��zע��i��a����3�ev
���p!�/��?e���F�<o�ئ�J���ȊR=/�Y������!3�]���2{$���kt�2"�el���������VP-��d�2�%W����T0*��&6|�i�ex˖ф�S�y�����wNN��lj�M�[2�5�\���[�қs����9V��N�dpKKu���W�����ddi�����Ԫ�\1^T��`]���k4P;�~�8Vb
A3OB͛�	�<�AMU<b�e�� 0���4�KٴC�eZo*p�Ϯ�C���
��S��qHkW�	�S���@@"/h�F[��M!���c��$f5W�:�8v(�9ݍ	�zP���+̔VUb���>�ްZ��>��G2��Mh�ꕁ}�3����f�W'@9����=~�\*�4�y�H��'�f��Sq%��Ɨ�|o�������>r�4�c��hJl��x߁�8�R�J�W�߶�p�?*�i:�Zp��Hq����ﾗ�������U�f���Q&�1��\��a��Y� :��ـ��z��
������oʕ-c�zI�O��VP"�3�y`$�zr�:)�`��<I�w�Dr�@�
o\+����ֲD��P�A����?3Un�{�X��,g���N���A/��>�aj�F����Jή�6̮���R��SO-�41�Fiw41U�:n.�,��n�~� �?�f����,���Q^�a.���^�>E\�MV�t�C�E-���)�iӻ���I�M��N�+jG*�8Y\�W{m~��ySܩ�ߙ�����9[�����!��f��%��WAٚ��~q�kZ�[��A� ��P`�M3$��֒�4/���h�f�����o@e��1T�y#�lw�[ժ��ڰ*���To�Ş���%.v�dr}��W��(��x�]F������L�B �c�c�5��ۮ�J'&T�v�1������jE�MBRX�PN�)
�	G.��� |�ʈ\1���kh���w D!GA�j�<�D�	�uG�s����bþ�K���V����	+�'dˌ%SoI"J����8��IhW˚��B7
áB�΢xE
~�3�$<��	ӝ��EF�}S����5�|CĭUՅ�QW*�Z+�����j� F=�(�JeW��eF���xw��(p
kW�Pa1^.g�j^<l��)�B6i��+�(�f����'��������v �,�ȍSm���ߺA��g�{ŏ��яn
̵|�����}́L�L�ley؋���*�3mD�k�V�1sX�o钬���5}rF�,���J8IEy�Q۪��Vy�4&���F"E�Y�H(#�.oəD��'�$]f!����T��
�	�1;O���/J��FCB8v��q�c'�7�V�*���NL�A��ìKA9QGM�~A�e_WyL�y�Mg<[��F
����q�-L0SHq��59!{�U�ӧ���B�,��9��������Z�B,,C]�Z��E�0����t
�A�7/Ľ���mr�*ʡ��񃬉>��^Q����F����#�\J�P�/La�W�ǊvA�S�`=ci��u��Gj�{��/ fg�g.^��+D?S�Re8��� ڞ[�����9�
�����5��y���,GL��Z��_�W3��{?E�6$|��I�R�C���_�����֢[�T���e��Z:-�iT�^d�-� ���K��=N $�p�$X^i�����߇�;A5����s�SSN@�n�/�+8W��?�N���;B�×��9��ec�S���ڢ�&ϝ����6(�5K���ܬ�|y��ˡ�8��b?4LY\�-bx���ףc��ǝ�%�tC/�ɲFQz�����o9� �$h�͌��*���0ZO��lu��Z�R,*��)?	���7F�U�kqn}�<�$|hi��H �:q��] ��G�篆���>��]��߫�O70&G�������r�p5]���ħ��M�)�Z���GfKR�q�Oe�&M��^6Ĕ�[�x	
<��C��2ОbV�G�qؽt�Oj����������K�y*��_��b�/����D�ʹ
Z��滊�<��������n�j�j@ϩl��OU;���������%*jf��F�<4���>�b.�(oʄ(pI���OB3���!����H�M��������� 4u�� ㈪����(z�Ao}�=S��ӫ���ҿ9e;��� 5�*w����Qh��b�D��u~cp��2�:�;�������t�^����3�U,�2�?uӴ��-�qɠ2�C�U�]?�S��g)�p�����T6</X����d�hF@^`��_�7��+sʫ��WWJ������
��z^h�ZBse�''�'�2*��,(u�
Nm&y1����Ǉw�B� ��a�@�3�I"fDB�
U���fΤY�Ƞ�6Ű�M����qbY���YZy*?�s�{O��b^�x� "�R#��w�뺅ɶ�*"�&m�H���{ �|�˱�;�X���3�?�ٺ{Ƭºu�?%r'�Fi~�E7�&i�z��9m���i:��V���'a���#��%Q�V���U�񆨏k�;CђlԂbD�"`G��O� N�c����/=��9������`��q�s�qB�X��-�����ߩ��(!HA�?R����%����p\�3�w �´�?u}�r,DF7[uB�D�2
"�ŧ����&O������z���i��7��]�BdP�E�D�K{��sboC�3( �5�@�g�J���Tri`���o"�. a��Ҷy�E����;0M���Ѧ,��mr���T��~^�U�]�*4��u%x֐T���R�B�3p�B �p,Ge0P����2 pl}�#A��"�l��î�~�X!�*v�0akW�>�!�X�������+�2+�͋���]u�k��X${�}<�~��_e��v^Bٷ ��
ZU���=#˟`vA�h;_���X���Y���D?��QAr@^W�����}
�-��_P��h�1/1�Y�$ ���PQ�����
��s�e)�e��-��"�����~�.�z�]`��=�qƋ� �c{���ÐWl�X:,g9��������ʉ�c�!�-�G;`�QQE!v/�)������ظ�$��+:)}W��F->"��R�����/gTPR'�(����B2q��z�'&����@�)��Qj�I������*\�K�	h��skuo�s�d:G{�`1�(
��E/��� l,�b�zB��Y�P},��8{�ѵ'���Vꂲ�M+�*�攇x�
�q�ҦVՍ���i��m��(#�?:!����nA��j��Q�W�����l���E�ݒ��͢W4�	#�1���e�pa�Έ��-��Ye�@NTyi �½m��s^v2��<&��R��aWJy�z����r&2��p��J���Z�u�YsL�6_�Hۜ ��T�.*RF�8�w�E%`	h�"e^o(��s�H�Yr��&u�м�� ړl��ɋ�7J����ܶ������K���Ԡ�� �\���.��Efk�^he:��Q��V��۫k�3�����%��J}{�b*YZ�:�x�#�
����nן��Y(y3|r��W�ւ���>�GS�I��F�Yul$`D�?�-}��������:��݇6}���A��'�/�T"1S�����,S,�뜱���4�XeH*���� !�o���6*�~���>6���m���ƚ�1I��y��3��U,;e�A��#�������.�c� ���
Vx���畯�	JҠF�d	u�@
�V���b�v��D+��yĘ!��!������6���?!O���.�I���d�V$�?n�p�}� �(>��c�OUyJ�VA���|����^.�@��!�@�$[	Yj�^!7P4]�Z�i[��5��]���9�^����� �U�9(W��ڋ]CeUv%Ŋ`�%-n��Q�4�������'H;��KE���Ȕ�n���x2O���|��Y���۫���b�'#�9ݪ?<<kv�*���V ��;�}Z������zRzPUA�JC1�}��PCh!�W��:l�ػ�za=�$���Zo=��x�Ѱ���<��eU }��0��k`�U�p�2I5!�3F��7r�H`��/_6�dz�y|
[֬#w�^��I&,����DA�7�<�q$�h�$�X�W������(�I��=R]��yMkr�)t͟U�=��+[%����<%E�S�N2��o�q�\���|�&�| c��;�\
�q�S�6D�����- �I���{��t�5�W���+�r1xP����U� G��kpڧ3���T)���LOL��oiu��MJ+�25������eM�����������:J�s�wp�1[#�\O��b�c�X��0�3��ި��0���h	.�?D~^�m$�����zI8�����s��%����O|ӢR�e�#�<�.Q,]�n�d��7����dBA�C#%��-D�Bs�8 >[hF� !l�~���)��3#up����]HH����1����b ���H�Y Xq�+m�=��W>�x����8,���zȣ�`���x=�r���ũ�Em���Y�6Q�>��_b��O4���e��3D�^���Rz�w�ϥ�tS� ���'I�2(�4t�3R�p�+���1~{�&em��?����*ƾXX�C�*�D_�J�&
ͷ�W����B^$!uqPe��s�����q������m��$GX��yi�3���i�%Is�h�o/ �+DT��P}���Jd���� �"��ǉۨ�_�h퓯z��.�(��M�G�ފ�'�+8km�y	<(9�_�n�|Jb!ɍ����@�f�tY�>� �ZF=6���D������t;;��ö���֘:�C������0��U��'�<l����a� X�U�lf��p}M?�bu�wsS�D���x�3
)a7�K�r&���<V\nd��8Dci1|i���GCo�M�*r d�w2�q|�!��g{0�)���X���:��@�s��0j�}��?@M6�5�-��+��X�H�W5�U��9���nP��o���Z��+�v�m�kd�:����<�#&�b��l�q��j�awq��dsk.��75Dۂ.J���sY]7V�ֵ!�y��뉥�k�!�/'s�x��HT��lb���y���O �=��{�r�#@K�W�G�"��k��UW���ϖom����a$��C3Hӻnq����b�
�5b�9Br��OUY���G ��J�Dy5���Y��Н=7�VMw7bkn�f0"9����`����#߶��.[~1�i��_�6n���?������>
�ߊ�f���&؂��O{��]SF�?ϳ�5.���/\�$�cg�58VD�pg��vdx��$�p��̐3�F�@����](!0��?��Xs���ݐ�_�Y$�(��1 ���}
3D1��<���j��37&ɑR&E �F�$)�����H��m]% �Y�MS�[s�S�-}~)�h�)N"W�J�Z��:s&��}x��;_W��[�{�2�7�1�,�ERP<
��~�:��$�!��{���|0�$���M�ƆĐd�Onu�x�%B���ܝ�[��+�93��T�ʟ����)�+�@��w�3��U�&��K}�M���f<�Y��0��ƅ�F��|
Zj1"���x2��������E�Y�a��Z�e��~^/���C�����ȤR�ͧ�&!�ї�����!U@2Y��!ɝ��&�:�]f~��Q&j���d4]�H�:�{a1[;�����m�;E;:}ف�9�K�t�:�k���`� �f�~�0A��VS?%�V�3�VM����!�����q��-fx��uOEV�YUR�һ��81.���2�Ǥ�m>���t�,4~%Ԏ�V�ui����VV%��Q���qo#l��������"�o���V�qK���7˪�����ݔ��-���좄�<�X���h�u�aW��4a3Z����kS�X,v�O����nL�Z��{!g{��^���MeZ���[ �(C��J�Tt')�>%�|{3�� �q�3z��uَQ"'��z�U�+s0��(w����c�hi�<S�`������-��ax�\'�V�:�����bbᶅt1f�!��?-��l���u�ۧ���4���f(�/���gMd?�����7���@�h C�!�w���;��mz���u��02��[*�QK�!g㸣��Iw�nޤ2�0�s#w��Z![����T��4����c-u:�P�#�����v����NI��hs[��K��x����s�W��C-�����4�-D�*�O���e��U���u~�n�ߦ�GKM�o�B`q�+��*��,H��1M�jZQǳͱ�G�/��Rf�"�������>}��Ȍ�|w�?�L@�"0.$&Ǻ*n�-��LB��cF��hƶ,�m���"�d{m5�qCJ��0����	0�;=��}���Z��?J�I��U׉#�v<i+ՓV��+�L�w���Ru�Q=�q(5����4���Ʈ���.�R*ɨǪ�l��B<cD����+�49S_�$�ع�+��&���\ci�"JT�A��*k��ζY� ��a1Ю}@����1�[��=���4�H�Z<���e�'�vT�b����tJ���2��KA�� a
���<r)W�q��	Q=^��%L�>���v��l��x��$��Dj�ޒJ�=��\o�N�*F��0q��	�&������/$�m�����V�;�3�������0ޱ(�$�h~�|�Y]�PU;��O)�<���pp���Ś�ʱx%z�^���&��;�L���V�]�d������G��q)9�����W�� kHH79mp�hv���-��n�N��}����R՜�_CxWO�WE�;�h��Eq��~�N�Wraz�ߙ�vo!�x鬉6��
�t�Y��6����Z�T�o�)�8:�
�U����q�Sf�%�d�(ܟ��>������#�!Y�3���=�]��8��i�:��Om�D�ݡ�����am2��i��������s�r��*+\��=��_�Y��n�0�=��"쵅��?P@���1j�@��9?����[���:���3C0�	�}Zo ��EK�U�퉇;���2��LI��h���	|:��#�~�M��("�!cg$��}�|q?�#��$_��}<Y
�<��#x忡�)Xyz=	F/g�$�B�߭�{�j�bsmv�4�8�+�"\ ��#���#����1�,�+(IpWSw~�L��J�؋���h\�B�")�V�@�_T)Ng)됎)�p���{��Z���[2�)0����g�s�
Ǵ	�E�@�<�#��!H�E9|r ���5GJ��U�r�.'���罧�lq)E��)�����.K 6��'������N�q���i�����(�?A�p�DR�`�B)ײ!��KY.0QJT{���&x�G[��]��LJ�uC3<a$?2�:��nbcZF���q��p�/:X͘cHi�RK[��eA!�����J���~��΅k1�Zoo�D�f�7�F�@1�mh��}�Bȸ�����n�`O�����IC(���Ԧ5WO�-���/z�
ߴ\
=%>��i��G#��aV�EzR6+ߡ��TBn�F��|1(��l߀��(�-�T��J��f�<��V�}9�x��C^�S�����::���Ws-�7��V�c��ʰ1؟joUr�f�0=<|X�ݣ��d卿(��/����oV!}��u��Z']*�LvqEm�3��/��A-	�-x�X���R�f�;]&��&#HsB��"���(�D��@xV�[�i�䱖aԃ5)���_r�T�q���H7���;=�����fK?x�������#c��Z��!��XS��k�����yB?1�dN�v�+lq��.��o����VT;�%�.=U�dER��kA����F�fo@�X�Ъ7t����I�����(l�{��0�h��zwZ2B5�k�7��N6��yk��}�Ҏ$��R�̯+>���D�����yqI�EQ�$V�������x���Rmm+��/��.����Œ��․2j`u�"Ѣ9ud�Td�!����K��x�F�;��h��G�uN,�0�ڟ
]�%�eM�7>��	���T]pD�#H�gs�8os5��Z��6�zؓ�FԊ�Tl��\��0^iV{W2��!��}�b���
���aкEv�m�0dj��3��7]���\/�2/���3�R �nW��ڝ#	/�#��o^��8����K�&�(�èiA��qڂw;0Y�#*h+>n�o��ZA�Tr��h�xaʧ�~�VU4���
9x�Þ3��˝�T�GK*�Bli� 9x���(�5�Mr쵗���N��I�\~��Z�=LO&��sN���'��$8c�Q8	;�!�!����.D�ա��$���r;�S7���l�*�3q�|���5����鋷]�<*G=GH^����d���k��EJ�z�I +� �ͬ�7�\�:�|v~H�N�`p���� |��E[�Z��~ٜ	�@�˂�_�否��ˆmj�xn� �*��v���ͧH��*�@K��\>���-����$5zv�w�*�+4
Ԓ�6��_I~�jX�9���
�F���-�a�h�z�]La��n\b%��]�JӶ� ����c�ʄ�j��.�r�M�	m�`c:��'�>��;�˜{Kl�B��~Z	�f&���Ǜ'�q&��{���ݽ��ز�>�c+9��U�F�A��.`e�J�����U�;���
yY|`T���@���q��q��K���DF~�1�cZ�G0L1^�S9"����v���,��8�Q�����t<�c���T�o,	$�{@%4�?`�4k��� ⻒�D;��A1"!�X���q~sқT�S�F����Z��I/+�Fx3+�����/��ʥd�#a�QZ5I,>�Y8%�錚u*��*��ޞ�t_�ڹfOT3񴇁m�h�
@y}��]ayG��W��n�j�������D@���H���9�.��u�������#fZ����"�F��,�;��W�ȸ�L��c7Y.=����^���z�����O0x7�6������=�*�?,�uJ�>� ��B�"�&��Q�7>�t'��"��c�U��t���+�x7�8���7k@�C��)�������sK�5 ��7��7�$�<��W�I�JXp����ނ�hxG��I�l�w0)�_[�bPd%�^�EƖPiQS4���JQZkE��|w�������0(�B�o�"�2bSA����	č �
<=�3�=�Ί/;�hɜ����era}�0#�&�`���Wj���������x���"�㙇���Y̢9�y*�n��~R���_3��Ս�"�1w~��8h
���I
�+_�[�ݝP-Ne��Ǭ#3B�����͒��Q�~��A^�s=��VT��`�쭗j/ݣc�d�!w����<�n_(��et���Un�>:������M�FZZ�h�U=�����ư�6I g��+�ר<|_P���He�����[�[u�"V�b~8�8rf|����K��a�����ꮀ�� S�Gq�0FP9�r�"0��P�"C��%�5d2&Fy*s�'ez3�!�x�]�QY�Wn���f�A]Ũ�H�$�v}*[��������lh�tmz��k��^A������ǥP������aK�8J!�R�m�.Aq���2c��';��`M��T�c�'m�o!J�t@6����$���n�a(�d8Gm0���:Q�{ӎRTd(�C�-Zg��3F�gD��0���i�8		�f4Gɗ��7� m��7��\������c�(�_(.�e���(�%k�)�#A�8U�tO�X�I�c2�+�J[w��K�Z;�c�l���E�u��M��`��
���4$�2�$U�b�h��	a���fC�#����Z�Ƙ��~�2x�6(d��O��>��n�	:�H�|��i�k�T��a�ěv4�ϞB��F���.Q�E -Y�E��-{�;=��h�eJ�~77(�Q(����@AT�^[��@<��W����^>pA�����5��.X��1+�G"j204��yt�g�{|wê$���ږ������۶�o�j�¼ڞNY�Wk6#Z�p<"������I���N�5��
L*�E"��v=�����^�.Z��qOE�*�ف-W�	X���-��9�qV�|�&����h�7%�O	Q��6�,�A탷���R�� 2KHU�)Z1����!�}����	&Y�L
��ŝ�D������>mk��ٔ�Q�L0�)��h��
7>�k�׀�}�����Ț�|�b�H��1��ې��Q��gW�~u�����\Y�>A��}AaFSy��&�����p/���2]&��H��&�x�O�$$v�Q�7�{_�E���Ϳ���sA�)�j�ݕ}T�5���qb5UH�d��H��5�&�"
܂#�Ɨ쬅��:vV_�͆QxԸEPζ�R�	����~sm�gPG�um�J/��JAC}?�צ*�q]��y->�8$	ED�R���	]=©ى�U���+���G��P;��D/-��ڛ�z�P�L^��2<>l:l�M9�j�'Y[s����x�;ܹ1�0(��N�
)�= (��̋:�"֌o���7�8fˋ)ZeK�Y�s�.��� M���HPNv�y����򿦼E���QƟ�E�l�%sf��P�S!C�g�CP�g��`Y*���8k�֧V�n�,�p̵Kq��|e���d
I��{
��tL\[*�+�/zw7�VdP�+���9���9��uj��$K�K�`�X#o�^'��<��h�4D_9��ϐ(�#�&�j��L�� ����7HE+4,sӃ}�N�8�L�2�"i-e�:� ���u�HăU八��xu[��$&z��H�ړZ?�X�9f��1���+�����5J&��K�4zZ<Ƚ��?��g���5s@�6�kK� ��P
�VQ?R��a�����b�U��Ta�Q\��Ny������W�L���KP#�b�L!Gm�{��+E�-![�����к��FzFu�<���
y��dտ�vn�)��@����uϳ���������+(S^B\@���f{��ۣ@C	jK��)�A�v����u�iCK"�PJ[h����,M��)�T�f�40��Fk�v�N?��ٱ�b�HY�b2�o�v���ȉ���ӣV�\S��z� E�ǀ��D��`�͉��Vۤ�I3�B�͚W׆hA�o�eH��
��+���*�]R5q �`����Kծkg.zQ�L�l�ߩj.���(�Pĉ��FஸøL}(�sX����Eإ�����f�dX�������^��Z�]=)� �^��79��d��[�Zٵ���'��`�4��I'%��֧i��D�@h薥�ؠX�k��XoR�Zp�s6�w񄡕G#�JD�,�J�,?7>������q�E�h$�&�k��+Bմ9ϩ<5 7�_J���h��@#��H|ѝ\��5H����]�57Tc^6 �
/Kܣ��}u���w�ؚ?�W�����Ҥ�l~�y�R�"�[�k�2����ChL��>R4����g�O�!��J��=vϤ�g���j�T���il�U�=]i�\�<Z�+[+D�8�ndz(5��鮟���P'��Nj��ͧ�H�%��]&�=�}̴��F��y�v/�-��%;�WK�,_ǿ�N�c�92�qY���9��k���4eז�!m "�.24z �+�$��n��>,q��"�ir�.����Ł)���&��i�/�՝��ՂAn%��[��"�K L���Hg���3�?��@}�gu�0�1��޸��٦"U?׷b˫R%0���E�v�����K	|+@{XV����畤�q��*��T�Fl��N�ɹ���9�)�����
W��~	lm;�f�1>��Mj���W5UvѶ��&���
w�����Y�O�Xz�v�f�JtՖs�g(O���x����s�ǻ|İG�G��|�	]��"����y�ф�Eg�5�������xocM��=�?��r��1������j��3rxGg�q�cŋ"z�8;{�2��F�v0钔45@����TW��q�����O��O �Dr�`4��\�?�����ak��ɗ߃��aif孈&T���#���M��<}�l�����z{S�����{����y�h�
Ҧ�o�I.Z������}0De%�_����)0�#����oA��b����{��g~��;�l25_v�߽�o�9\�Nb�K/<�7NlTĦy��x��W��[ZYjS����uL�7�z�	2��s�u�U�e�{��E�>	V`n~_�%y�P;���q`�tN�x���tb�*CO������I��Xg_	�1�:o��U���3'&~�S����t��9��Rȝ�i��`�A�ݚ����m�6��Sր"�:�:��*(?I�2���uH}�o����6t���&� ��͇��ϡ�de�a\�<%#F��k�З/
9p� ��m�z[�Rd�R�n)��!p��顨#������u�����N��TK�A����_�SVH�(�;e_�XA�=�R������IbH��46�vj���K�͍	�G�������~���a=/X�M��n�����a�?�>��w%_gU�\��:�������w)�3G�PAp��xyb�6�?�~n3��*Ϟ����`��38������i�+��a��eu����Q4���:�N�LM�YPKh�ēo��Y0�@0�pă[�$l8y�=���L���������t+n�i���C�Z8rN"s��O��~e��߾�x���'՜[1�f�p`�$�)���o�n�us���OjӤ�0��K/k�m,m��7�	O���E���%�s���;T��T��^��ܝ~����J���]������;y��g�UV�� P�����/�k�b<��s����7�v��0���OM�`e��y�ڀ��R�	�	��@��1UZt�tf�+���
������.��?M"�3��S,�K�O�4a���'Į�v9�!ʋϟĵ婧�G9!Go�{|0��t�,=�f%�D���2Ӗ�+�簦�S�[j�V������-A�����|�\�rvW�+|�Ƈ��/��xQ��7�O��:e�u������������o;l��y���6����g��4	a ��^����ǸSͫ�yۄƛ�����{��LN����-�ykeX������`(��I>NچsO��"^ް�s������P�r��h7}��(��t)J#���=��;�Z�p�-�CU>AZ%�u).<|���3�;��<�U�G"����^6���bлl�RZ&��l�h��6��IG�X\4����7��䉗�����-�C�Ke�#�*��M��v�U}T]�N.Y��-��y���l�pQ���q���f��r!�i!4"��]�B��KX9j0
z�؀dmЃ�uM?�%�CC���p��Wj=�^��/~�1���A����ͯ��� T\�O��9tv�*bm�
9w>K������E�.����8�J��ɦ�[~cˀ�{C��Ӵ���-�k�����Vؖ��kRJY(�@�,�y�=���`9�N �ƃ�"�Ʌ�����ʆClM��Wb�Y�N��!��|r��d�g���e�{��H���W�c��Y5Dx"�r��X ��-ιM�7W����.�[&8�Ӊb�{a�s�x�23�D��$n��vA}�oݚ]\�X�g��k��U�o��!έ��a�2x���67��:H��8`���vYy�4o��: �\U�mĳ��ݷ��Ԅ
�o<���UVU�'�'%$e0	ͅ���d�	4��Мc�<U��@#�4�ն~8D�*
>� S��v9�<�7��K6"e�I��]����^d�y����'[_��׶�,=���|��I��8�2L���nb����M7Vb�Ŷ
_X��M�������lLC����3��@
�=��#\�)���V�3��?�i�^�U7��������|+^�c�����!�$�'��JP��Ms�}�ջ؉�-�v���[�Ԃ~:O��}<��=E�`V�u`�Xa�V�K"m8�����k�,�Ѻ���6 <��7V�x����
09@���
�w�꘣9&��I�B�!��kR��:,���b��_Í�/���D��������QH�����E
R�����-3��8����q��AtN������Z��(�w�3\�g$r+���罯.�������@�(T�(*�%�����Sᡩ�ķŌ�Z�i��@Ł�[4Q&�b���HgH���z��ɹ�����s(�е�yp�MϢ��]q�k�� �/.�m��K&�����a
Ӹ���<
˲��`oS����y{2b}?��$����O��|���a��}����3ګcB�X�=�ڗ�񖌡'hQX�#�4���X|���v&����.eWWZXu��uvT9:�k@�M�i{���cK��9e��}��rT�>�5�O��J��f��<U�{�0�g3d[Y���q=q�&u��p"������6휁�>
�"�5j���`� ���'1�/��>��$UR]�pc����Edʣ:fï�����;Y�e�aq�4�����$T2���?#�� mGB�W�ah��P��8��Т)� 댩J�#���\�#��+P�#Ӓ�XUgA&�3��"�b9"���"��؜T�ᛪ��DٞS�y>��ZS}ݫ����������4��t�>Dv7�i��R5*vB�dS�����m�@�#�%��I�b"R���@�Hr"un���1��`�NyN �M8�j��$�� 2n ;��gѧ\�
����C)��W�Va�+��]$XH߰`I���J���4$3�ZS�Z�t���.�&���p�b�o�`��My�����bbV���!#�<'��6�I�&׉U�����qۇeJ��P��Hub�U� в�ؗ!�e�2�`φ��4�v����$Md���U�q��E��%��%V�4�a-H�I�O�\��U���]�jٳ`����@.�ù|H��������dj��`�GZ��%-3�hᢖw�_m��-`��+��q�J���|�[Td
�}���1e��3a�jd��O�>���E�?(�vb|������*���w���gJJ�T�;8�nҀ��g���w���9��!��Pҝ�O�m
z�'΍�Jb`�yzPnJ�&�����u��I0-�����T�΃�#}h��N�2C��j��	��Z�-D�M-Bm�ak���{�9L����w�Q'�W���1��L���k�\(h�#+%����DgU����4=�&����S��	/7��-� F�ie���ڣ�i��4�~�A�L#{��i�����TV�h�2H���,�>"_5#�e];�>�}�A��y��6}絗_i�#�m?��Ѩ��G./��VW�݊��01�!��r�p�̸�E7����D� yxU�*Y.�C���1u�R8�2���K��D�.��g+p�}��	8�E���|UwՆ+KD~�p���֑��h��6�@h�r�"��|%���rZb�԰���;{��5Bm�����gA8%CC!w����Y���Mxgj�<��������i4���ӭ���Gy(t�P*���K��.@�g�+(��I���ix���{�b���n+���'
�>��K�6�K��ٝʅǶ v KV���3��Q���_]��䶍g���@&|�Q;|��U�B��z<�'o�Z1TrQ?��ܧzs��i��P��+�u�@�4�K��њ����_��s�3m� N'��s^�WP��,e���6��k)@���x��E��ޖ���mR��!�	��FG�*�m~K�L6���Rc��&�Ǻb՘�>�ҿ�Lb�0-o]�\k,�}�ܒ�O�o7��(���q� �vv�}�:A�E���SS�%I��{����3?�:��o��n���4�E�R�;���]bO�`�XSCX��q�d��T�.�Y��{'!/%�ŐI�g2WQ���@�x�,S���'��zn���8�
����@-sR��q�K�w��N����,��0����l�#��A�?�̋l�M��@��e��E�
[���d����jp~q��*�!ɋH��"����O�o��Y���
���u�uX����(޿I���5Ew�%�yRk�;I��i~�����&U"�C����j)�>��Q��8��\�ܒ/�f�jyk!��/� �V,��\6�Z�_BIˍ�0k�
O�4n�#�Ę
BA��^ȕ�򨌱�2ˈf�� a�3�?櫃�M�C�hӝA�"�)׽>P���\.���/w&�9���WP2S,^co��=����Ļ�Ɨ��<e ܦ3�]{�Ä���#ٿNG�%J\�Q�wb���`^�C�}ۖ�"=t{���D�h�C��V@M̈́_t|i���a��.�+�l��Ҧ9e&�%��t�\~���]Ty.l_%��]� � ��A�b\3\^I��O����k�"�e^pQc0��F�Օ*��GjxS��Wr��\� UA��eb�k�E�W� a�Hi�ȑyk�@�8��.K�gd�I�L�>�o 7�����}�.BH��XV��Ks�z�a�[IOh'J��{�e�<�G�#�<�>}��?�M�\�@���3cגx��չm���OBUR��o�bB�W��4��Z��Cb�lwT�&B��i#��J�_��V�(���>g�K�^q���%��{y��&�o���=��TR�n	�T��G}p-}K�r8��*g�T��ލ���4��(l-��pxA휷+�9���"�=�_�`�p�vpf�1+"�dsf�M^Z�mG�����Z&����Ļ�q������N�c����Gj;���3Kg������l$�r����y���+iM6�}�A��W���F��?�ILX�`�n9�Bf�y��mk�C����4���jU;��;��i=-N��y�c-5p
���;	̼�\��X?ȁ��l���.�K p�ZH�SCp��^n=��M6����]�ČH�Q�"#�+}u��o�8X����u;���q1���"Ic�8�`!���E-~N�����h�q�"�ՓLY�'/�?1w��$����}�$�r���2	*�?f(�ʤx��r��J
�ұ��n͚�a����	��������~tz�Ϥ�,�'V��a	����������2��$��x��{v��E���_��T����
�Ǥg���h�t��_��K�ʩK'�E�]�gY(�L�=i�$-�6usD�q>�TGM�:�z!w��=w!��x3�R�V�c��r���K�b�9����% �-&s�d�	�15aw)����!�Cf/�q������1@H���
YJ̀�Z�8��87���YvX�1c`jd���nP֪O����1�+HύZ�i�p��nnH9�l������H��1�t���vc�%��"{,n��ǣ��T�߶�Ո�h� O1Y40�u�dN�2��ZpD�l�����hz�_
�>��#�r�����m��j��P����uS�^���?$�$Q�o���Y��|~lE;��ˇ�墥����}
äZ���X�%Un�^~-L(i���O�����4�J�c��Q��N�Ƌ@�,����O �IV��V���5Btǧ��ШEl��}����9
g݌�����~e��:�!�sa��$=�Oiʊ�s �_���R�8��/�������y#����3X��YQh����^�T|�o�$�TI�:u��Წ������N���7��=�<��;,b��c����i~Ym8<3�>bü@��?ͬ��79��s_�w����7�(~���~����7LB�RB���x<�#fw.�x�fk�k2>>̐�Ĺ���� ��?�'���
%z�R���>A��@�`+q��Dx��w��
~�/�H�o���d)br�@�1-�c��x2�P��$��s;Mz��-�A�{���W�$`��Y'I~fF8��,x�6�㓋�{�����C�+C$K8:(B��>��!'�x8�&.H!`U�0��q�0�Jr�9j�H�R�=0��!7ƫP�B�}�T��W�!�&�p|6���h���:�7����C��A`.�j�|���C]��O�ᗪ���~, i33�����!�����U�s�:�4*���3	�6���>�dR=�>]�D崈ʬ&�Q`���iG�]\N��ja�\*Dp"�!m}����RF�B;(�<L��i�e��f3�8��x��ļG`3��iC1�7�(	�N��	p� ��2�yJ�؍�ˮ��f�/�E���ȮО�T ��&�v��å��`A�ڒ��7�y̒�B�ڒ>��D��¶x�ŲBY��,{x�Q�B����zR�oS�]%u^M�����[n�&��E'W����DgP����}}�0���w��tah�A��0�⁨�BO�!����O�FLTLC6��G�����`���Zsi1|�,� � �Npb"\}�F��m.C|�15FI�2:2����c�Ҳx�d�n��x�j���B֗]QI�	��Y�1�>#��R%�
�q+{,��S0���F�꧚�;�]ںtڨ�O��l�I��C��84�`'y���>�|׶D�T���;���ՂA�Vh�Q ��w����@�����_��V$�%�|&�O���A��H(/�	 ��
�]��V�'��(<6� r �7;� Ř�Ə��ť7-Ψ�fi��OC��
���S����晫@#�6�@�Z�
@�n!�=�Y��1
�蕏$����5��[ΰ_T���o�(uPjW+Y���C�3�'��a�Vqu�X����s)�&�۪���s��a�ґ��vٸ�%����y��
=垒:Ak�E��m�T���p�.���F��o��z��ۆM����0��p"��5�~o� M5��؞z��/Xyj�j�f���4g:�Ep�M��p�'A�[=���^�N���^�RB�F�}���%+('��Y"�����+���ʼ�A�������O��=�(��*!@�"�"�L��G=r!��
���O*�݋��bL�!��Wj��� �	���<��m�s&2�}�4�3�O[�98/�N���Q�j�<m�P�Grfͤ�|uɘL����ZC4�ruP�[�	���y�)�3�U3	dF/��wܮ���i�Vv-%v�n:�I���Θu�T�BB�Z�OCG�cJ�l`I�<)V[$)�~��V>�j��l�k��i�ґ��2�QN�b~8�$~(�����S��1�@�� 9���L�2,rMQ��	�6���P"��C��Ց�B<цJ�f"�&�NWWLcEˊZ1��2f)B6������U�F�f��<�̢:��Ӯ&wѨlЖ�j,i�i�vX�U҉x�e�h�F��t��]�"'��߽�y�A�M��D~�[��D�~���g��M��5J:<�������u��(~�y���P=�*a-&m?e��Ug̩��9q=���>���VrŶ+�./�̃���_5��R
���>&4t}�����rcM����E!����J,�?��������%�g�~���������4�����#������9t��t�V�J�峱(�����R���7����9	��ܓ�ya�b\���W�s������P(q�8�l��ah�C�1�h��ř����;��~uc��1m�R�?�VYm���2�+���X�ѝ��}*��v��Z��[�⩋�V%z������V�4-a�q��Ng�@��q��S7c�&�l���bj����4l˭���Z�43�c7J&֪J���	����Ͷ�k�!|�N�M�-�\sg�
�^��B5�/Gu{�=ŗ����ԑ�Y�^��~xL��?Iш�7-�X��B�Br�V\�l{ׁ���`/��4.m g+~Ȼ�~������_�"]E{��|&0>��]���.�ڄ����:}�)^gO����:N��Yj�)(��	A�`;-�������y��K`�g�ncY���sg�{�=L�~E%[�����/ܿ��0�j�Z.�����ƭK ��ȫ�W>v
O�V��eMfD�u�(4�:�[0tͮ�M�aS�Q�����(r�"y l����Y+��#��h��܉,~�#���
��x�?���dm�L;�/�-���ڼ���b���rPr��u9V������JP��Z�\_VQ�zEq�iѦ�f��>g�#�Uȓ��A�c���̓*}Rt�m�M�jB�n� ��z�1�#���-	�?ʡ:��%*_����(�.��W��N�y�+r-�W}�ޢn�s2:�$	8��5HP�����涥���	�q;�wu��@�� ���'p9����OZ�[���?d�9�K�@ݪI����$���$��H��xJ�XL�r�n��||�s�3�{#h����CH���1�#�{��Y���N�r����Y�{7KG�E��(  ��f���A_0���~&�"U�B�&m�2Sh�����P�-�oO��cʫMn�#��tc�>�)O���Y8���|+ϑ۵���Z/42-`���V�|�"���O`<r
dX5�>��@�ܫ��v~�#ۼ5 ���P�88�����
	�làhp�|���
�Ю�>/XL���n@��(�DW&O����څɝ��<zdT�N������Tٹv�DA.�m�q�3�DoA�C��<�5���A��z`���
(�ΥS��'dTQ���S YB����d��?�de�#lC���u�(��4 ~���9�Mf�ټ��Y�,���[ԦD��V�R.&����>��^t�"�Y��ޢ[=�x�?�˼�$��"v�&���^䨴$}Ͼãt�QDY�.W�aTpi)���%�E�:W��8�%� �}�a-���f��σ��X J���U��qre ����ˀhʅ{�\�羣����H����Kq��EH��x$�O�5��Y�s��p�h�e�O��L�����j7�2�gl�˻��8��2*>֗�45��Ѯ\6j�����q\�a��x�sq�]'�e�
0���fh�	U%�L�y9�C}���b�����<����={m������lq���E3Q<Y�C`K�nA��"��� }n&t�]��3��x�� N�Y�����%���\8G ;��'����Uޯ�D_"bwD�w/td�#�x����:_8����ʋe`��P���.�s��i7n�x�Z�Ay�"����I4�0do������y��F�r���.����Z��խ��^�9���LΠ�{�f���8�X�j�\�?��� 
��*�$����hB�o���T/Z1R���p�+3iMJgiz1Ưa��ߊ��6`E��)M�Թm����E���A�K�埻��}���zk�1�U_G�%�.�8]��2�3:�:���ڄ��:���}䶚:EE�3������}�VjF�nm���[MW�d>0��W�Dp�qigsx��]�"2i0�̕=ٙ��F�UH>���ro6�S�KNe1�Ҝ��K��[�e���1kbN[�l�t�����U2I��d�QRR�~���w�������G̠�}}#�\�>/�m�޶�[�I���)��l�ֶP��y���鱁a���c�Du������s�5��ߛ�M��'ψL��\��mt�>�Q*l����r
�x�V�SUq)��u�9"e.�_��.���7�«��R�,Қ�]rO��s�E\�4�Ct�������
ǊpeA#ȹ���7ãԤg,��˗{��H��^�;1�)����q�Ju������l�B4�v�1�t��3�v{岿���F�|s9S�� W���>K����|���=�����rS>[�z���������\9�ۆ̀���������Fq�ܦ�Y��o��	�ѳ8>0�YKD����c��7�.7N�������w�Zv�֍�iR,�*�Q��)��|�>@M#�AY$JlmY�|ō]a�zL\����Qe�3��������+���O}FeO� ��a�[M���O�~T*��vY��%zX&�E\�"-�����`��F�K�~}+$1��y�f�3�j�g����eH ��V��N�W��ե�s�]�O������ht:�&��u#{zs�X����du���O˧�#��H�*�E�t��Q�r��Zq6��T})Q�_/���D�R�C�!QoC��u�8n��Z��D�<��H�<=�n�LB�lHN��V�hZ��ƾ7�U�� ���0p�w9������xkmW��1lZ�b�<�9���E~	���܄p�ui�]���3K�8LH\�>}=�|h��u��17	������� ���n%�&�����)Ğ{�9�Q����g-���^��y�ԩ���T�Fg�ϱ�[r�k44��	������d�:��a4��˭�yـ{�����!�耘��*�L	m������*��є���gA3�oUܝ�+�`WY�I��iR�񽪰cq^S_|:5�3C{)R��2!��q���N�r�J��g�z|n �GVH�y���ܪ�,���f%��Dr8��[͐(���WJX��e�W��PX��d~�c)�ޟV"��2�݀K��Y\����I�����2�k�&;�r6�O=t��RS���G�]^B}`��oP-�������\v�?��������~���雚�؜���ݒoR� *����B�����w ÆJ��@/���H\�ʫ	U3Kr�K�����){s|�5�2ӭ�}���!��#K�)C�2�	��+��١t�d}� ��ʅ�s���)��#WM�/c����x����)b�6����A�8M3���I���UgQ bY��
v��I�R�2�qF'8&�G�m�i�I�-��X���C�f���Ee��?j:�L6��D��i����| !̄�Ta��u-<A���`���e���e� ������ܷ���)w��<m�,��>��HNO|�����"��l��M�4"��-��F7G*��Y{�&t`���XGB��k�Z$�����;��z���"�P��2̺�gHo�$O��\3�@dU���^��*V����AW���'!@�U`e�����)U*W�~7O�a��s7���\��q+�.Bj�[]�?�I���@::��%��W#0W;c�1�.5^Uy�Qӊ �S]K�A��I@O ��|��2�T�!�Z����ӡ Kf^�u`������y����I(7�N���1h��P�#Ʋ��2�Q��]���Ý���^�.O5��hFI�sn[�qW���\L�=,8��������WUɮP9�D~�n���*h��H,��-#/��r�z����Qi���+�ㄱ��W+ID�#Ι��ɏա�n��9�R8Y�����k��$8�XP D��[�-\Nu�+D��K9�b��!H_J��F�P�0��.8�S%v�.AME@�֯JC_B��zѳ4�5�a�^��MQ8�|��9\�CE?�������=W�T뛘���㙍w��$ "^�K@�!���6e}R�ҘJ.�޹j��S�K���0�1y��L�Dwԍ&�z�m�Mu�$�G��&�����*!�>[������=΁�f&B��,+A&˨NPGw��ܻ��i�a�]3y�t�|��rN�먅e�:sȞ(�7#X2��tS^�A L
i��u5���G�1.Bx��{�v]
[+���?�Ri�X*�U.�l-gZ�!�=�!p���T>��nҮ�=�U��A���P&q/Ng�6ƀ���ˮ���K:t�|d�ekǩ�&�,P$���#�xR$�@��>�V5J����PD1��J����_o�$,FP���))��.j�n�hEGpq���u��P~�����PVhF��wFX�,��=<ԨD>e	"�sl�b���'��<����!~�����0~�@x������*��َO�W �~�ꞩ�՚������>��t�+ZW�K�u�:ԥ���Dį�����z��oˀ�I'�1��P�%�j�ʼZb��8�кw^��A���)6N���=������p�W�:}��Y��M�Y��@���1�[^x���ꌻ�JE4�zo�G�r+A���b�0�9��_���ޱ�&m8�!Mc����)��B�)��M�����Qi5�vͩ��b8��Sb�ص����8M?�
	��Q����9�\�ɴpEw<�G�ږ� ۯ���q~Z�_����Ci��m4�kro�E�DB�oh^�q�8`�Z�fp�%K@����V]0��גa?L�@������s��d��o�`&��(�T���;S����??u�O4_r�dqBg�šN�b�t�tW~�*3�̜�^z^d�1),I�"��G��/I��&�%�p�O�G�B��٢���o
�r}@X$Y¬�Ztx&�N݌_DFj���:�:=��#6F��jǅ�qf�s���4��珡!Glr�H~	��ւۭ������!��#n��MIn�~����t/]���_d�e��7^�v����}�6A��s�������?�]�S5C�鼛=��9)oV�F[gڞ�6a����?��s42>me*@��
��{��a���"�2��~���o��
�
o��uTp�N[T� S|w�mQ{�;���B���H6+�������K ��Kֹa̯��L��Y�?�����������+�f�< }�hϝ�{�2ò.�j��5�y5�����.B�0���Q]���\������4(�W!��*��f���v!�f�#Tk�&�^O�8�6R��3<q��QP���-�2�}rN���c�t]Bm�BY8���0[����:����
�+�}�T��W~��OX�ʷ��G:d.�KA��o$�ץ�Xv�݊ђ�k�\���H_�uÌy8y��$F�Oa�e�D��5��z����F���w�	���|n���Tm-X}7O/��p�I��Ә-�D@�����֣~�e��%7^S�v�$��b�:Y�LC���b�.�m�<xwc#��JZ{�E{V���j�����Akd��g���d�n�[<0ݬI�Bh&�;�p(�u�]�~п�?���r"�4c�3��P �~�`,���˶*���J}Q��ߐ��^�7�`_D|x��08�L&�o�3�sC���a~�Z���7�K��h��5ge*�&4�T�@ܹ
@Bȥt��o���b;�;%���R�E;Ϙ���f� z�묱WԌ/����\R
��O6^Lw�)��CVO���j�^0��Q?�Zf=���n��4�2-p�{,�Ӻ�)E@�,~>����3�k�w��4-�M�#ik|OGq�̸�%b�� ?9!J5��kX�(��FԞ%	������Y���x��DP�'j$B�C�fb�4tuoma7e���ͽ6<���FA3���V#��)�1���$ƓR�3MҞ/ϭ��me��J���G&�l�!B����Tê�E
v\��h���DK�r���k��[R�odBD"�B��Vww�߃rUy��[��ڋ�5��^E�a���i.f��?!WQ>~�S����'st�lHTo�~��f�r�JY�D	wM\�W	Hpv���0G"quS�2��(���C��ZJ{�]�zl�*��?B(�J�6��b޷�Ԓ��l��֛>U�=#�iB���a�O#��]:�Ԫ�>��ˡ�Œ������q:�� �+�����hI% j��Y�͡��A<cŨ���a�yż�꟟J� \�b>m�r�ϕ鉊O��FQ�5��T��NH�`��b6��
g���3AY(��'Z�ǻW����x�� ���z>0Ūxx0j�E�ژ��l��4~�4I�fh���/h�&a�!�zD)R��jc�ye��Cmeh������G���b�^'=ǀ��?��Nm�VLe':yHU�����ՙ;��ޠet�	��q�1����Acɜ|�^��B�~_f�]|� ��@�?B���B��`sD.����� ���� �c����DU�]t9�.1��UL��tC����|Nփ
k3�����	Al��������[�n7�'���kEO*!4N�x�\��]}k�-�%k�_�����7K��X�_SdB{��7V��P���!yK^�qC�Op+�����Y;��	�*��3�h����~j�Qe�hxi�Uَ(�3$��<���䩠9�o��L
BM��$�%V�����x��#E��;J�j�r��d��#@-�h�+_��k��ς|�MD���GÓw�Q�ǋwא�~���z����r *��oҜ�w�G��������` {B��|7�f��ҕY�<�0-O�̳�[�{��E*!���1,�>��/��(m��u5�& �Ǔ�A⃽7X>)�c�����$VW��q�E����g��+�\O'�{�dqL��q��A^����-^������(]����k� >�*&�}V�-�Y��J}z��S��i-̈>Z������xê�S�Q��F��;�r5�բ|	�.��WO�K�U����JﺖNC����|���Is�P��E�g�V߃��ͱd�sb�M�b]'P�. �;�6���tp �rq���='�<�J�Yv�D�]�j�1�_�)�nb��h�ZiuBÞ�s���ݖ~�E/�ȧ��g���S6�ǹ�%��u��q�b�����Zmy���JV/�z0�:��.zȺ��W�}�-����J	_���ٖ�ߚH����[����b��O�| ��Hb����?4t�C"�������-���Cp7S�qZB�{����x�������f|_��Ȱ�n+���ʈ�@�/Hg?̋6��&�I�3�����U�O��P�D8�(!�O�"E>�:ep:��Ե����ń�֯����c�_+�XY�_W8����ξ�(�{��؏�-}gռ�u�7g
'�;�@-���$j�b�WK�=3�+����]�
u�M�UK>�S�<�A�<H��t����X�ݳNX��T]JVx�;�2�A܂].s���ջW�,c���1�>&P'\�U��2�s>��G"$n
���g�}.�M��h��q7��'�'*�W.~�l�!ntf�v�a��,K�G�ō�����g�9r�),cd�# o���s'�5�\u:+�n�t|k���&'u��yW��a	
K��#u�#�
��۱��b�b"��Z��B1���WUJ�>s<�j/���+SN#�~<��3=�̀l��5�̺���P�NqE��ܐ!�0�bL��3��h��~�f��Ɖ�u�����ƋC� v8���-����Y}�ݕte�^ج�D��Z�=q��P=�y}�Yjq�����	f��b�ջ�ԟ�� ���YK�ջ ���>=3g� �Zd�\��k����H��³I(�p.h?<�泄�Ѳ���6F}֒�cmŌ�����2E�1�*���,��HE����O_EMlˎ��5�S.��R,FB@�'�8���P����vџY�{��fu�@e}J��xܾ1� wr~ n�$Y��xv�y���H�a�8-�Бdi�=�p\P��ESFnE�@����H@�(L��5_����"b�|���Փ?�K�o�>��]A�p?����	p���H�&>\��k�/fj�Umh���d����Bb�"������Qu�8(`X��y`� >e����zX�����h?d��}�����>�+kwW�Z'`oW"�`e}����ܬ ]b�͙��F(�
uN�L1�4��ο��������S(9���9iIffؘ���8}�����' K�k�"a�
C�����dϝYNnR��1v����D�����,��}��4�d�P$��s�]�2��+~�5�o��|a9�ӓ~����m�]��g���򮸹��dYu��i�ˌ�q�9������O������@^ΔJ�I>�Q��v��}��'� �r2�mǽ-�G ��A#�z�i_r�b��"� C��S�w@����5B�@J��\p�W7KS�O�-��D]���Y���fy;N��#.љ��(xn�Ӑ; u��~D� {�d#=y�b���l+��!��S sX[#Y'Mo{�N��f!gBK����DPD���;��u�	_PH H�ecF�����y��p�|k�y����E�R����Ln(�I�8��tN��N���a�9�Z��]ug����X`�K��z��%v�8
5Z���?3�]��	+Bu������$P��Zv�}`9����i�1�W�����47*��Hᓵ&W]Rd]%��2��?�(�[��B�0���c����D�'�j�Mld���PgVf���9�F�`=��Ju��G#�H�E���6 m)3�1���#��[_�^п)��+o9��`��O��m!� y��t�vDP�F�OA1��]�3x\�$y_���J��5R��њ��oll�zix^<8�)���'�W���W&.	o�0]!->��T���!�������������[\'M��eQ�c�fXV�d��!�ZPɰ<Z���[�A
[�oe��62d3���^�B �1�dG���L�߳�ϼ�x�l�O����]2�
~I���zj���5��0�m�ϒa3�5��p�8�҉3�
{r�xHeUy�qq%�ʆV��jya�u6��,v��1^�j��C�2}9�C>4~�^?WY��>�����f��#)�{��>R�Gpe�A��V�MorCg���̵��R|�$�R�ܧ,eٔW"��F��ɓ~�gd��q�ט���)(鲍�ӕ}�����3�~&�Ns� K#������qI�w�D�L�����l�+ֆ��Fhp����A�Ӱ�������?�
{���g���7�kJ0��oOC���>�-��憊)�|��'�D̘ΖrY�����z�ΎTq8��?GxUp<�Ǽ)��Lě�ZM��_����������C��	=x5C@���KR��"�I���h�7n%bs���56L��z�9���Q�N�Λ�-P[~Kȵ��x��*�C0"�x�#��^e-}}N��fOָ<z�_�δlI�?р�D�,<=����}w���z���<ep���r>b�	ˣ<ڙ[hl�N�)����eҷdXo�]�����C��w5�)c~u����'�@�T� 7�0�u=>����+���k$�Z��ݿ��i��!�0����_0�9��q.^�O����^9t&�y��rja�w;�om�ܯ�����B�i��(
 �3�%'���c�ln*~���h����1Eb�'_�77��=#���ǟ�}�_6ꀃ�	 ���2�jES�'��v�G�坖.��$w����ݕ�D��w��(��f�mA��ݲ� �PH����R���iw�k�r/��5L�k�
�cQ�"֧߀�dZ[�S�0�����7E
�Cg�(��Ru8y�9|xݔ[yZ�[�n0���)�)�p�WrƗ̽�o���6�;�!t2[�S��+rZ�P³A�/�+NG1ur�^�GG�`~:"�&�}d�*4y[���z(B��N�:�)��Q�d�8���fX��PB+h=�V��	v.����`��_'�s |�����Rs�p�n@���M>[�������g�z�,�pd͹�D|r��k���a�i��	R<�l\�ڃ)���'�t�B��1A�K�-5��Cd$IfĽ{�Z9��z0�ȟ��uφ���e�a�^3��R�KJfV��ܟ=s�f��Ã6Q%e���u ��36��
��VR��k�Q�@�	{ AV}b	�$8]�r=�f��6N����(�j1�va9f�/x~�Eɦ6d&F��Vڝh���i#'�m��]���s;���g�[�u�8�ho%.*��p���M�z3.�!z�u4.�{�q�#�t1D*�+�!jfOp��3�Y���C�v{P��8�����Ƅ~X~A��w����%&�k�m'Ӥv���Hz���4�7��=e��4�`��h�?�U!��yH�;?	�X�ׂ��,�ŏ�8�
LG��%�:
����e��̨l��Z�6���?�ՀvE-�e��� *96� t�i�
D���S�K��k#11���2bh��������k`{�'I���[-a�|{ߋ��h)�=�B�!���	��ME��O�Wә�P�C'K�Nz� k:���_у�-6$c�a��?���EH�_]t_�Ea[��y/U�$���h_=- �$G����d�����KP���R�H�,�8x��ϸԜ���
�b���8�������}9���҅!�?�P�o��z2)�����-�Ѥ�<7���j�<�K$�����F*ub�Z���|�71��QX_e	;�y�>}[���R0��L7&��~:�P@[�XБ��;C�%eC�&�揓-Z�(X��V��͢���osJ!k@FDZ^c�if'�4{8ņ���ģ�S� e}A����^��&Uc�_Z<d�s4���DzH/��W�k4E���)��y��&sм�22V�QrR�u�6v
����gEuͮ��V+w��?MzT�U.h��q�k[C�$4�[�כG��=�/�8�c9j���e�x�~�!�-��O�����q��8��AZ�
%� �qG���g���0����g[EJ��U���0F�;�u�n'����&���t-|g�ޅ�hv�}NJ(�t�{�&��o�q��{ċ�q�E1������`,b�Db�-o����x���Ϩ4��x��g�&�_��'CohƞDI�Z�Ѡ��B�?e�oD������f�����qQE��@gI8��O_`�0�P��mƌ>D�p5x�h��y�Z�E��_*V�:�ݒh�}�b@��l��0�!�Y�c��*JcQ�����i]�
n���Cɰ��gH�-mҹ��L�#�MDXl,��;ȶF�B]�u]
�Ka�b+@̘�����I�n`m׆�S]ɞ���1�7@ �G8��L�Sx6�d���f�����K�Ӽ+j��&0]�M�*�.A���{e�%`^UUS.��)���q6ٹA��||� P�d�eRwً��^�{���y���Ïw���n�;�\T���:�I�y�3y-���@j��n��|#�H��K�7���MRե¨��Y���8����kGT鋃���ܶ�$�^N�5VvO�l�HT<�����ݚȎOĽ�,�q_�14�.��sxZn%J�L=+Ǒ^�5绋p����S�z���z�0�Z��,�Y=�m��lhN�HR�m��6��S5[j��J-`��YĮ�sь�&"@�0H��C��Z S� ��bH�ż�.��u��5x" ]���aA�m�B��\�|��95���{O?�`l���,r�g_�$�n��87�B�o��`ez������Q.��NN��ku�t{j��?���$h-��o��2q�R���x~���A ����q��R�(}߮�	!��K�6S#���:K*��g��k���-%�c�,��
��9t �)���cB���z��K�V��@qh���:���Z+�1��\6�i�S�柼��͆P{)a���u���`3fVk����쐏U+g��j�fB"��<����0F��4��Wߖȕ6� �2�	�Y.��>�zh6=�i�Bvי^�Hц:p�Y�ހ�ݶ1�:�`�
�
Ċ�i��e�}{W�6��3����i�O��!n.U���ؤ����w���-�$��T�3�{`�b�&�Q�p�k>쮉쟅��##$���Ц@�f���=��
��-G`���gd��Ge.e�P���]�M2S��~4C�f�-���镁��>u�q�[Wb4~�4�r&�I�&��#n�|���"�F���m�L����a�3v�L��7>Xh�0�>5A��1w�����P�)^$pꘀsފpB_�[`�}�r��ϩ�#cl5���#՘�%b�I6yG��s����n"���y�h��"/<V}d�t��T�f�V�7fǃ�A;�
��C���.fB0�䟱�T�I�^C���(���o��2<��,�n�Aа�S#���C� ;��X1���z�V6]���\�.�Q��8 ��0_�
�ǥu�Ʈt�;�p�lf�N�'WL����_ŋ�q������X�j5}J�j��6-��#%�����)p��H�Q��~(�i�9��b��( �*��¥"#zvtq��)/�&o�-�Ϻ2_�}�;�/�Sכ��'��ܔO��(K�B@Q�����mH0�g�f�S��Ɍ5B�~fG�Xz�Y����A�b �����PU�:��.��ږ#S�M"���Jo�M�#~I����zE�	w��ϳs��	��?.���皯4M�3 *%;�W?w�O,���~dJ�m�E��E�Z)^����Hi�a"�ȓ,!vV|(:މ���*+2���s�l{c�� �`��<�j]��M{W��9��"�eO�*/���@ރB�<YL�$��nm{�5�	#0��"H7*���1Н������M� 
���򱼿�{��X[/�e˨)�_.ٵ������3f���w7�t6��_�q�Mc�M$P�q*�s*쮈���nൂp���Ovx�m��'Ѡ����i9�_ں����D��ɢt˸�a#Db�>Rꇞ�2�z��3��?(�B�4h&���q6���JN��@>vËϥn�N��<N�������e\�6�7������ed���`Ѧ��F�	(������6��&�D�rOxTR��"�&p�g�݊���K�V����\)�GS0$�4=���i�v�	���&��(.*��	��#�Gĩ�k���&
�c15b$���4=V�B�d���WY����Soc���/�U��[b&_�o{���/��|���In�;�F�o:J�����M�6\<.
�UhT-��Is�fq����<�8�o��`!j�59�Z?b��V�Z4���`�f�����k����ĥ�	ŕ�:�B Ҟ��ӓ�k�(3
�~���6Y�^���'~�'o7.q��c����Sl�쟕=����+�����SB�E������?���>-�3��?뜴3J*��dT�U�m%��H_S�ܼy�62�܃�!�@�̎��O�@�dd��.S\�ong��n��>T:�EGH��뙸9�P���uF�`�Ue�n�&�}��5�OdDWx#g��ܦ[?4�GO��} 
�˕-�͐��^A�o���z�Y������N����͕G�,B��k��o�Cd����ءb ,N^�|��٫v��V���_�GE~�)_P��V\ �Qwx���\K��#�������0��~�ը����=�Sv��� Ke~.S�"mLC�a���݌p+9����^Ɣ�A�}D�k�����j2�wS�m��T��op�0�H'V'�i��~4����Ի6
00D
�?�rlu�10��#�<XN���+T�l�e}��_�H�3��ҦD�0��w�M|�������L��@���~j�耨�Pܸ��z�ӛ�w-Ss�����_����%��ۼ[%�ݧ�c<,�F�,p��,�N3Tum|����si���ת�m������?(�j;N����#c;SJ�}��O�hZ�/�9z<���]��W{�����x'	�*Q�B	�_dt���1D(�R���4�"`0�7mJ���"��*I[�B��`>m��?x��� �{G�Wϯ�����h��X �_�_�q䥎w�>$#� MZ���a����=�q�+��~#ds��P�N"�� ��������;p��ѭtJ� �9��!����Aឲӷp||l��N���?�ڸ
%ҞP�������fg��$����v����q y�|EAM"���ɏR�"[��@�m�г�J�J^�qkͰ��.���)���0��j:�͞��A�28b��uQ/��9T��6h%���K>���ϕ�8Y����V%C��+窆p_���xBꩋ}G��8�+(�����A��[$uw�R:}wYY?D%^m|�qj����S7��˗�A���c�ȏ��
���~���F[���K�Ê�g��;q�~�-|����>B��*tJ��vP4�����P�fOiP5��}O���9g#� H9��15�3���c��e�����adzH�1��b�d��k�{�A���	\��MP��bȡ��������ons����<B�c��ŷ����c"��P(c�s�2�_?9��o׳"D��)/������٤h�u2!�ONn���"�j>�[����3^�OpQ��o�g|U�h��CWl�E����^F�Q��Zo���
��DF8��Ձ�+���	�ܽ������r�n���a{�Ĥ��,�����x��r���1?�Z��Ww�b#/l�y
��^G���&�(�ro�?�uߦC�bB�����.��?��k��l��q0�L��C�����L�NC���8?r|x \�;f��{_�r ,���phF8Y�MN�vo���rk���M���S��p0@�v�_ F�-H�^�2��mU��-E�XGC���^�����en�E�2����d��?II���	E�:S�e���jʾ�<(A��نȉ�T��p2�~a�-jx������}�$�����z.[��hu�һn�|R"��bԕ���H��+���J�ҷ�W��t�"[�y�J5 �oE�ȋ�ӯ|f�4�~0λ����ÙY���aQ�s<�����.I�[v��gߎB�mM�w�w�H^�rRO�<���^���{�~<��t���9��5�'�4��E�.��<�,��.!s�H��]���ֲ�t.�T������B�CAq�]��j��x���zv� �cnC0����˿��9J��/0A&8+���Y�R��\����*`��ZLr�댽n���k}c�5���D{L��l|�I Y?;�AN��#��H�s��W �/�?yU4����<2�sI��3�����DL�I�b��3�s���W�"�m{�����/��������SRg�wiŨN�5����k�\�lHKlV��^�\�����;�o���bg��:M�_�1�U(��*�\�zĴ㛝��]���BQx��O_�	��Xt��(�\�iz���5�l��T��͒�	@t4�`�A���m3�h��y�gz� �,�k �\��+U��Ӗb���.	�z_d��cc�p��Ln��q���t9���HJ� ���ĩ$(� 3c�W��:J�� �� �����E�ń�
pɔj�y�,�>����Ȝ�l�&�S��9��*͌\����������_uy,�;��Le��|{-5 �\���u��)��&Wy2Ӌ�/-�*4}휥F�
@������K�����L�"�f�p�,*z��x5��d9v�´�&.�zE�X����]Р�7�;+��H�,K�b͟z:�ׂ��"u�Pl�Ei�î��~�^�^lL悞���g%�4一����kn� �z�n��ӹ�j�>X?��f���E���� q��iJ�ߺ� �h���H�\���k���Fyt��߹k��NeOF�uh�>�'B}X�ɒ�A��� ���Γ�C�u��fr�����s�ZRt ���X�Ra�����|���DP�ސ�o����dW����.�
wH`�I�q��<�9��P�9�Qz�U�+P�ȉ�K�>e@В�*�Wn>OM�t�'*.5�DmEoa��K��4�}�E�1���F9�\$��@��������D'?�c�Ѫ�!?O��C�Kso_@�`��KdIt̯��4(�Zy�q[��\GKi�����5�k#��*���j%���N>���b���[;+e�̥_��x�G�*-��_Ѡ�&M�-8�*;{wk�UWZ�[��G	:��;:�uT�v��ڇ儴K��P=P��C4�b���$��� -��v-���M�1�kZ���ITh����
B��%=�l�%�z�x
o��`�t�[!`�Dnu`I�)�c��������*-'��q�Y��͢2~p}>k�[+�z��!�:侐uw!(5'�J�xR���!���g���j�����
���ׇC&H}�ǈ&�f�&�(n�U���s���F����HA�"J_�f(i�A%�e��O+5ui�#�T�uq~����*�Mt[�/��Eun��rv`{��觷�N��g$p%_ع8q��J�=���[4X3�)M4&"*h�ׁl��!����]f�v~��Bǵ�Ru��4u�{�g�ޖɛ�]v/3��������mI�Dz�	�kWK��UzZ��^1�S��MɊy�K��ʏ|f��Z?'^����q��N��i�3�b�z9��;�q��-�A�xƱ0�nX���s���q��׬\�U娝i�=��]�#4Hv)�cR�S�E�d���:�}�{H�����A�^o2�C��L��A$$�1|@(�Ҫ!S�r!*D1�j�+�/�:;��H�:��ʊ�Ҟ�D7��|�e�B:�YQΪpF~c�)�ؼ�!ӷᙦ^�8���\�����t���)��"�f$���v�uH���0�i+��:�e�k����<�� C���\�r�w���۩'H�sU�$3���;骀�$>G������Z�Q�}�|	��Т]��<�7��1��&��Iw-���k�!��٭ǄXby��s�e�6H�2=�m�x�M��	(�����վ��@}9��e�����s�A�!�.T�����ڹN��'������j�����I��V��1�N���Ȭ{�'���
1�R�lz�m&��dS�y�{'e,��4�ˑ�dZS��_V�!l�g>_�]�91%Yn��Qu�F�����Y��)a�E6%����&CjH�e�Fc!��']p�c�i��P�0YD-k\[k	>7�s�%Zi��:�y�U�Q�~�0���d(@?�R�
�
��:`Lf�ti���'��*&�u�r������o����z��+1�X���$���ԉ��B�L���oۣ4[�흙�1�Gi�J�3��L�6P��}ht`���D��E5���q������<'�Ʊ	�RʅQ��C���8��򺇛i^�Q;��ȯu����|e�����
��?lq+j�G;a���K�����Z

O�?�6��QJ����!s�57K>�HSkA�=R�o.�GDL-�0X b.�y[�s�WCÂ~�� �!��A���.ٚ����D,$�����Zp�B\~hN�����G�>l�R��#8-Z�;�C�3�
�Ds@F̒�	a��~�t4�v�Oƭ#��`�T�c]�ҳ�}�OGi8�3@�g �J(�>s5��g�]�{}I0��`��>�B�dFr�aE*~t�<-mϳH-�7��{�JDyvۤ��7ٷ����ϸ'��xgBL\B��}z+Ꟛ��H��R(y_�����#yD]v$1ѻ�Z�/CI|��5z{Z9E�F���ĒNwbC�%�Y�1��Ͻ���+������.�xZ�1y?d��u�S}�^dU�Ln&�yv��+�YH��4j54��MU^shb�]R�֢��s��ͬ����RGH2���F�'�m�^?/y�uTs�X��D��gc� 0J>>�����^ܪI�ǅQ���i���:�A,�&~���@�G���l\�]r�<)-��Rp��F��-�����?����>^o�W�ںZq�˰�*�ZO �ID��kz�N��[����7�W�g�8���u9�J��&j�:Zy>	�6Ad�:��գA�ԹV'��v�&����[�%��C�-^�x1P�4��^�>���M!�nD�$�sg��QxQ�`������i��" Lr*�1KG�1�Q��9�7c��\�,�~�)r�����?�Hp�$o���&)��o�ַ�ˤVW�]I���9-�&ط���s�� ������F�R��5���Nh��>^�_ۛ���mH����0!1k�cz�4M�2+S������D��>���J�K#Ol}����מ'N�Z�_��Py3�����~"�N�⛗,X	�D����G�Ư�P�2�uſ�z���H��t���I8��9yn��>*8v�A���k�#����O�ߓ����w\ġ:�fу)�R��m\� i�5���񢇊��F���FŚ�Ur�5�	+i����պ���6���[~b���aEZ:�+�t�N<�Ġ�TF^��E�	A-�(��_܃pDu� �U�_C�e��P�<�vgO��f[��S\i_zZ��9i^�Q�9ߴ^��h�l��gZovg�%�:7����U�.�����=�V�)+W��4�(=]q>��x����{^��kT�:�=kp�KК�j{�;Ï����	�"���!��%�%g�ٝi/�'l���7
��!p>D<�
H; ����w@e89��8����ˎc�* M�����P�Ʈ��9�l�/4�ڋ3;+��.���3���@?�C�杼�F��p��-��&f �]�i$O��&V.QV�"�t����L���6`:�B-vѢ<�(Hn ��������<�A�%�?���.7��(<����M�`�j�_t%������0~���$W-'�(��F�Z(��w��O0���X������j�� ,r�e���	�	���[��Y�﨔�l��`:�^��Ƕ2�h<{�R�:&A*��܇��K�|r\��ca���0�h����tz
%n|��@�s�2]ڳ�1��4O�%lT휷^Ыvf�����oN��jw�RԒϨIM���B�q`N?[X{�TZ� ���ZģP+Ɨ�Ț��5*���-��0)NHp �m/�:y;�6�"K`����.t����*��
�Z�g-�ELή8�e�I���{�.����e��.�'��~rB����5�,�H��<��78a�C�'�����eu[���T v�@L'(7O&�A��}������+"4�F�7��lh1��#��n��e�)��!�#�����U3
�%ok s������@ٷ�bY�����?��z���=��O�ޥ�~����+��1>r>ɂ��? ̆Y0�0����}(�	ʙ��3�=��A�	b��R���<	*)<w@΁�>`R)����i���kn
��̆�9䑞���7�w�L��O ��W|)���B��yf*���}�MQ�f�\)���������f4y�eC��";LMtK��twޟ
>ޘ#D`��<��M��!��Tf�����}��E��B����<^��r��0���_��h��χz���1��k.���uS[��JA���W�Y��L����:c"�Vm����L��`1���u�3# ��]ʑ���ѭE�a�3q�13��yX�H�T }c�
���Y�"�g�n�n&���&"�Z��i-��_K_Զy�1{�Vb�J�s�ɰ�0��NL�i}{��@@���j�	����
`�`E��b��S7�i���\n[��/_S���a�)�8F�c_�o�)췔���6^�TS�T�XX:j��b�f�J�B����m�Aa-���>���= �:}U�~V� _ذΒeo>��q�Fk�XZ��k֬�g�e�������X}�q��_�n�8�R����0J�k�\�7�@�w���+�\�ܢn�vQ�ѭ-&Ι�2��1j����Z!�9Ϯ�KH.���r�L���;_���!$񓴂qÁK)��FeL%ɯ�f��$�%(hI����:x:�B�����	�,}��֕�����T7a�?ck�n{����`�,d�����$4I�E²ԃ��(�^�c��� P���+J���t�� /@�G�,kn�U�;�A��D�>�k�XR����v�&����jS��n��`���:�rڏ֫d&-6��"i}�˖ҡ�Y5�-��
0��<\��(a����>��Y�v��][n�&���xվ[H�}���q�0�R�O:��k��5E�w����g��/�/��+8�O�!bڕs=�[��P�D�������f7b��;�Ͳ٢#�|0�~�a��V��U*�1�Z'�hc�P���B�d��avLD��:D�����mJ�H��30@+�<�H��Ӊ[4�V��U@��Xr#�'J����.92�Vd�87�9�e�;�b�q4F�Φ��Ȃ,qbp�R�8F��D��ƌ���R�`�[�۠�Ng����xd/W�¤$�`��\t˥����n��d�ю	p�n���ܞr���"���fI����ӊ�{͌�����lVd<H��� ��ؓJrz�	����ɖES���y�G�vćWҤ��HE$Eb���� ^GV�^�ؑ�>+x�xw�,�=�kZ����=�BC�<w��<d�����Da�k�
�|2� CZˉv}�^��soQ���=(�3�Q�`�ъ�̲L1A�HM�So�"�P�X��$�+����Qn>cT��X�u-�z��3���F1��L��N�w����ʪJa)���qJ� �8Lz.�L���ꗻw�d�X�s,ne�k��C��`l1ZU`�l��#Y�7�*2z�� *�Z���W�"��6�ay�)�f�
���F�>P|�g�]?y��v������w�N:ֈ5o�T^�>�+�ө�`a`��b�O�ɬij;���I��V��՞�%����#u�d[��&-u^5ő�8�a�x�a����i2����Ag`��h�ĥ�U	0�e��a#�X�a�-���w�x��; E���w�t��y�!b\m['J����
��H��G��} vw�ˬy�8�:�*�����@�Wnf�%�[:���>7/-@qݝ�5�J�4�����:��cg�D�6��X'��; ���-v�U�,)��ci��)�߻s�Wl��;�w\�&�za{8=$��5�Ҭ{2ɂ�W�q9�H��)�<R,���$QQ��V�{A?�Fҿ.��b$J�b,p}fl�-�A�g���u�7������xR|�uIL���9��]A��֗�	5�x�R�;O��h>�	q�!{�g��p�����(��Ż��3�_�m!&�$#V�Ev����o�V(�J^$v�Tx��g��B�X��e�[��ݱ�eDѠ�CPQ�gj�(~��r@g��Of{;w)g:|��$�`�r��!�{�@�׻�������jv���R�[K�nf��NG\�b����*���ٳ�FGBo�,-�E��!��t�2�?)��U�}��d����r�k�
�	��-:���k�$$m�Ll�����?}�ه�D�i�DMz�*���ۅ=�.!(KW�B�%���ɱ�JOV��.H�MH���:9�?i�O��n�8a�_7��K�UT�9O"���/��q�����ŬU"r'��Q����|�	�.HBa~�+��@u�����)�c(Hk*̤�x�$�28)w",gCODJ9�L�~,�fS��A��+�����k��� $�Nu��s���L�VT/�8��
CZ���k?z�ST �R=!}Y�g�q%����r�]��c�t+d���wU�$9�A��'�Ҙ{0L����q��xB��죚��F�+��E�4r9�Mz:�O�kK|D����/iQ+���|}�{���=����~r����6��
�v�;�>|�iSTߍ�̞�v���q�h��&
�ӛP�Q��t~#�wit�Rs��z\�~m����\�'�sK��|�r�Q�u_m2���[��}Q�Y6'��?�)Ӕ��`~��m�j��pYu7����=�g�u�-��YƑ������Y�0��.,�Кٵ0=TԕS� �8`��_?Y��u�gr�>�[0��M�����,�$�V�d��|�C���?e�Tw;5�2�Xԝz����������14.ZW���`�P
n��TP�WTEC����\UAx�� k0��ڮ�h��(������f`�TJ�)/f�>h���*�w���b`��,A�'q��h/Ȭ�h�=�5�����+%������4:y� �FUE4@��Q�|�i�a/��B�a+o�}#Ne�k���� ĩ�%.�Q{z)*>��)إ��W|�ȏ%�r��R	�e%B�A����_B�"�.jZ4k�J$�6&�\��md'��+�4�U!��g�o(��nc�F��6J��y��|EsE�-�J��OZz�_�� ���7��b��x"�p�M8�9���b�������!}�Wq"+LbB?��& 5�#��^��۵k�=45��T�q���)	D y��ۄ<x�-w�4��XQc^a�Qh�d�X0�$���D�\v+���b-��Rx(���y:�ǯٔbJ/U��;�����9�Fg��t���V%9A�w�Ž�k��A(�5\�p��X��70?@�`�u���s���Ύ݌�6�f��[�~�eƨ��Bc���F1(y9��w�m�I���]��M��7���[1U6G:D�|�9 �Tu&����	$3ُ������^��@��o�2F��C��d�̣
Z_\������1����js�u��X���wdv����i���a��z���.�"������J/�~X���@ؓ��>�ģvaȓ�W"~d�L$\5�:RSv홸2*dDak�;�js�g~K��N��u������SR��}��+U��c!���C�m�6K`��cO���3��$�<~���Y�
����������,n�R�� ��������nϵ�o���.`�ot��Ԏe�X[�:Tu�7%5lH��u3+�����T�����vGA����W\���Q>t��o������fYn����y].�圈�k�I���g�i����(��x�"������]�?sYs�����G�;��m�����x�`F-�$?�����Y�<a�����M$����]�0^�]T\ݵ���c�(��1�>S��x���[/0�x�Dai��Z��o�wNl��7�v�5Zr����k�`C|�E�ץ;�t�<�xh��H�����<�w(PX/>���h	�?�Ζ���$k���3�HͩC����FIA��~����3ա��JÂ��%�NZ+�~v~��6�D�+��NX�lr�8����G�X��C �P�����)H���:k���M�B@��|�����cZ4�ʉ�ъ��*@�U!nՈ�O_�N�� ������PIZ��:=Na&�N�Ȱ��2�c��ɫ��N��x�U�NY��B����~x]��l*?���DNa�������g��.�|���fݜ:`Ѣm�6�+V#濓B�O& ·�����}Dc:]�̝�������)��C8 ��#�;$9+Z/��z�}���:*%c��:�%kmt�� �'[����U�3o�����&O��*aN�iA$��{U�|����I_�'~[�<Rd~O��áb���:��8nU���j���\�FGVq0�"����Y��G����ђ��1���^��B��6�1����_�f��Wsl2Ծ�lKLE$0���C�1��0,Ig�����+��v�i�����c1l4��QM�y�Z7׼�@�(�>+�7]OAEc>�H����Nw�k]��m_��[�#�M/K(���6�k���� N8�AW�-�Y<���_bV�_%��u)��җ���ZC�}D/GU\˷m!K�NYF0u��qA}b�>��
�����zk+���#���i�����Q�=vE��&����@D޶z?'�U�TJ������k��i�L�a��#J�++H�ۼ�-ȽP>��3�����G#�ʮOZb�lD��&�s$��ߘ��� �hsiMh�ɀ2i�/o�x#
���v��a �c���7�UU�#�`T�i��5\��r4��!řP��^`�x�����˛Z��R�3�I�1{�x����� ��8�$Sp�ࠜg��ʼ閛V�T�F"�?�L�f�ϊ)`���%����>7��]mU�F\�3�`�zw>����)��*@6�fc�K;C]l(M�1w�.l/�B?>U�	���c!n�'��!����'�E&��3TfA��i�9է���&�՜d���<�����F�AƁ��*�+�~�k=`��jE�A�B�s�>�"�n|T��^'��`�C.��} g�s�N��v"dY�u��@�/;��������!��`�������8D��Ѱ	�B[՘(D�k=����]�n��İС�2��Y5�s�S�9�|u�z�*�X�768h�����U0���ΨD��ӵ�6�č6 �r�$��7'n3c�=y:;,#����L}��_�����$Yu�Bf�.e5L �a�%
��f�Uqq��(�?yk̵�m�� �J�B��d��+�Q�����e@���q���?��eV4��\e�}�7{iVΤ�-2��*��ޞ9��M��X�g-U���~4����F�҄�e�`0j_�c!�źK&չT�oی?~!����ު���٫���~/?�p�<�����5��8���3]�oh҄*Vgz�O�*�{!���yn,�[�����u�̄��ZA6f2����Ay�ˊ��/�#�1!�i)o0�9�h^���W:Z����˪�J/�=B���8�Y����Z�������׼G`b`�����dy�I��{�㸎�RdT��9�ĝ�R�q�!�U]�"�ک�f��ew���pHX�B!�0��:���~S������9��0U�p9��&TrP����C�9-�|��z�*1��f��oB�b��z
k>�R9�[����Rw�t�̀����n� p�
_z
����� N@ �j��k�5S�#wj�`O��~�l\�J�v�m�U>ZS<
��z�8\� W���4 ��-����5�y�}�(
�w)�"�6�Sچm��E�&���P�EBN"�3$��ڈ\���{�w�s�B)wn���C��V���ИM�<�e�:�0@�>A��5'�bw�8L��i�l��.yiL�@��:2a�@�y��������#�3ݣ�1�����S9 ��� ls|��a'�bq�`tMډ���<��G�:������l�6Vb"���-���M!U��%�ጧ���zi��=J���|�-,�A._B���R�ʵ#��jY�����P�8��M�d �m$������0�6�¥���7%8>�~3dRW�:�Ԓ�Hm�O���6�P����R��g�ψ,
���Aba��P�e=����4��VFg�5����h���(�Ynsi�赪�]����#3��<��Tٯ߇�i�_xÖة�+�33!�_�ڹf���(�4�ﭷ�/�����0��ּ�٠��w��&Q�pa����%����tJ�`����Y�y�Ʈ#�΂���{�$M>,�C}��pbzSΰ���g�S�����-sb,$*J�7o2PD�,��A�di����j;���|	:��n�~�{gr-���b����Y(��"��YK�Ϳ�B�������%돨�D�c��k��������c�j��ࢻ�s9s����JÉ��)��&-�hT�d�X�_��_��R��@d���k�Vr��A��V��C}��m�9#�����Zn�� �׌� ��.s�D�?�}}�C/B����a���^>� �V��z�v�M6Îc�:�NN	�'��x�l=}̏I�ŗɻÑ����7���OJF�����΂�2F!�
�(��[�*� (��ƴ�o���G�TŰF�(�hMG��/�wͅ#�(��z�͔}) ތ�8�����\��H��� 6s9�԰U�}���XIs����Wq�x\ibq���FRm�0 +����Y<�Ve���!W�s�	����g��=G)>�`Vj�
���1ޫ��y�K�43�A��P�o�5�t;ɷ������v�wZ�qM��ڤw��op�{�!*P����4��5�Ew1�#���a��}��R����m�i�	K�A�whU���G@�^Ѹ�Zӹ.��2o�L�C�.udq��Wc���o�����$����G:�lhL"kN#�4�
^��x`�R�Iٖ�u@GKӗ��C���86��	m"i.�㿡l��UG�:�,/���H?����D�D�6$t�Bc���cִ���ǿ`I%�EC��K��hl&wL,��` �vac9� M�ŻȪ?�F��=$�ٷ�5���ո��H��j�K&,��ÇQ�|�pv�W m$��7Q���SuS����|�R`r*����-c�N�'` �/��R/��{i��8/��cb�A�Q�m$"B��A��'�G�c�g��U��������t�G��O{�q�������-�����F�'�Q�:?���.���p;�*3���L2����P����N�yc��N��y�����ri���g@�a�!��[6��u'b����W�y����4��Pޙ9���ؘ	NT��Sf,Д!��\r;u�6Z������T�h1^2�r�H�� lnz��g2L
��@e���cXyn"�T,�T��L�I츁�Z���w���W�t.!�%m?ir(��(�����M�m���("��|��}��ứ��:@�����d,�/�BK�8�/�����?W-W��cBJ:m��/�C�&g9�U/����a*�^{Ì�^8�
G���$�T1�D�iP��I�^2I@�Y-4"�ǒ0B����&���A�5ڲڄ�$������^-n��{���2�r��_���+����ظ��[��ԯ��}fH3�\;���j�B[�x�J0d!,�M��:��x�W�u��T:,�W�B� F��w�`���-qAV�ŭq���l��ؽ2�]8%o����C�ۨ�A�b���ٳʴ�ngل�L�
������Rfa_ SN����d_E?��4�<�-�Dx��x��%|m;R�Ld�{/W�s~Uï�^������% Ǽ8nj��4�T3IUAPtc=�����e�Lp\�G�~�3�i����5 G�Ǡc.�Dd��T~�*��4�����������'u%�~�����R�����Ҳ1�������L�h���(Py�3�!}m��ds��|v�N~(��`2u ʸTqs��sp��q�i�r��ȧ��q���܄5A��dxet,���(���0�[�>Rɍ����J�xr^�[z7�2Eqf:�=���G:E?���_��,�!�jc�R��>a��efT�L�����NC{��G�=�-� `��e�F�8	=za2�T���E���,5s�"���^p��~�>�/�r�FQ����^嬫�y
_�e��B6%�3�������k��<���K[�g���'t�s�*>P���7	�mI?�0Iϲ(S���tM��	�����O�̠���7`��w�ͤ�9�CX��x�Q�$~�}V�7fm��7�a�_���w$kCpi#���lp[\�j����=gM�5�(�n��S��Y�!����z��g�9�M5w�+u���b�bı�E� A�$�A&gw}�o�g�t���je�^��χQ�d��l@����C�2�\��M]V�Dܻ�d���U&m
�V/�y�zԼ�!�$+�' "1�n9���Z�.�8i�C�{2���;)˗-g��!��{
�p��T�
)g��KHp`�L?e��g��^��\�0B�r�ϫ:���<�ħ�z�vj���N��C��o�I��]�ut�x:J*aY�^�#HE�2�c�ż��Ώ�s��Ŀ��Qa�P2�2�<p =�w�E6�0���)2F~Jh
��B�v�|n֌�����UT���e����(c�uo����)� ���%��֒��������؝�̸�U�ój=$�����v��%dŔ�d]���ە΋�r&�H�v������1n�ԑ�J�f����.  �?���L>�k�?=tym�%}/��}_��'�s���W��4�E	TB�Fb�=p�v&����:P2���������J&��2�1��#},�;��@�k@�t�lt�5��ZIu��j��CL�/�gw��JJ�Y8�>i5#��l���ݨ>� ��M�2�D�Q���P]x���ft[r��ċÐ�*����Lu'��0�Um�[�+\�h��}ޛS�B�Y*zXGK�JCaZג9wh�e����[�ߖ7���]k��`Kܞ�6���7qV���i�(C�y�J�Lzq�Ү��w�A��7�Wޕ"r��|�wЂ��W�����LՎ���_h=V>g�E�1[��B8	����ڧ��GLX����vcP��W�~��]`-�(�y�-342����lI�e��
KE�D����R!��ΰ�~f���!��Ocr���^��l�׶D.���=�0ˆk��)@�	Kv��4T��K����IJa�8�_9�5>��*r��r��8cJ�=0�S�A9�	�
y��'4Y���߃F����Ǿ;HXI��9Y���}����>��2��R@e�_iL�l�H!�G4�i!�
���N���nV�s�4����"_]�3�TR�P��LM�Hdrl�)��x�kQYnC�Uu�M��R�l�LL�-V�$��W��$ā�u��Sa@�l#EΖ�*e4vd��L=NI��e�S��@�s$�^A��aLV��`�z"zp����!F�hEh&��C���'Ow�&9i>�CH��l� ��<AZ���Q���޻֛�u�i@�U�-�E6$x�Z�@��\�d{�ok�
{T�I��lz2E:�"��a�4K����i���0ŵ�R�� Fu�2,��
�1�u�	T�}�;gЍ�H���{w�P��_k�+	J��/U���eL(HإI33��U�P+lM�u$M��`-?��9>;
-C7,_�s�B��m�JP�N������y�s�h}�����ҮơY�?�%�+5��UR�߾��L+�����"t�2i(It�r�e�k0�ϴ��j�m���sh�B�c�+ ��G��rJ
$����q��&��rm�}s)|b�w0��&�P����J*^��|b�]IUQ	�\aT;P'b��P�1��pRxI��G�!���9��c��5��gF����v+S�*X��ym��27{�l�_(ZT�ј��&��?X�#	ڄE���S�e{�����_0f�xu �o`�5c_)+5?�-/h0y�����}oef�gj�L�R�����������Y��۞�Fxj���S`{ĸ�@�a�N��(�D�lU�N�V���UM���ԛ�Z�b�!LyLZD��_�1�+i�.sbH_�l	П�o�ʯD�`1@_0�|aT�e+�!���Lc�g{K�s��#^�o:�xuP��߸��f�v��s�#��Fj�En�t��*;���r�e&5�gP��-}���B��	=k�ۆ�RIj�If���c �K�2����^����wr�a`���ʡ��Bύ-�4�8�I���H��9X(��6"�I��Irǜv�:�0�T[k	q?�r�iSg�D��py�Fl���+i)��(�5�VWR��4`̱�vQ�6�&����:�0x3g�W.z�E��H�.͌���dX��F��r����2����hm�1l� �&G��~)�l
��%����!	�Q����7n����ZG�t2vVCϗ7����e�@��gtp4��t	H7̫��6�b�~������:����3ҭb�73��if J�9 ����5��>cf4�-���H�;��l�T ��{V�`�G���?��̊��"G	k��c�lNp쯬��B�h�v����	C0����/x����xQ� �>z�!��UO��]�{�*3$>���mq%�d���5F����J��7(J�����?
)�^?J8�zRBe�5���b��wq�
��ϊ��s��8յC����.��a�ҳj��͹G���8�_�y�n�����`��Wc��X}����.�Ye�Oʫnk��S�x��f;O˘r@�� FG����?�Q՚95!ظ����R0�gO���f;'�Ft(�;>�x��
{���pEu�ƒ�
�88�� 	�������i3�D�4������2�rr� ��i�m���o�p9�:vZ#Ǚ������_ʶl>���ڮ�@�`�
�̺y
Z���O>���2��j�Å�T��<�P�ԅ{qa��3�]#g����|�OZ�zM�nU�<��e��"�|d��;�|2�	Q�H�`Ţ��ni�	K�OxX�ω����t��mZ��7+�O�:G����:q /S���\�+��dn�ց�#ۛ�Z��(���~�N�,Q�{щ4�X��z+G�ieMXC�����#�0�f���+�D����'���5���w.:zU�hvG��7-V-,CE�FG\!�/������TỲ��DdR-&���S4dy}w}���������F��S;A��m��A��5��B8�H�C|��~��%ʷM��;߁�'��,{��ޚU�
����q����,Êh�1�
=����O������D�#bm������ˀ�|sX�`���؆�£��<��dk�w�nE�u�� ������8"u��ď۾,s�&ǅ���O		�R�p�p ��Fv!>�B�9U�"����6��A��V\R'�K)^���mm�!�g���]�JH�6t�NgI��q�Nۊ�s;r���n�ef�C���0�uX�����Y��A�	���������)3�~�HV�8��~Y�@��}�%1:U��;��5;e�#��U�������-���V+�<�1@��ɼѭ�9�nH����@���lր�|\o*r�BX$��J�彆D	�V��H���e`�bM8�Q���R#���P�:�]!V�2(�[��m
:�Z���\��(j�M�� ���e�)��_�{�(>�n%`���ϊ��n��#�}��қ3�q��0��<��UE� ���!'SYg��l\B����T�Dܑs��E�OOW�D�TC3��ʪ�S��=��<|�oC�.����Vb���&�~5$�bE܄��ҭ�E��p�M�������넮䷧`��V�˂���5N��XS;�rm'k]ܡ� ���i�z��& _{�춶a{�7"~x�C{��!�qk�J����̻����-���3�	�=A�!ʌ��P���	@������*~�~����T�<���]A.�!�pK��T��C��ZA�_���Ug��9T�3����ŪHM��J���v`��P_p�$D�*y�ƽ�R�n�^��	�}Hh�`+S�K ������s �R�D����ez㻯۝�m���#M97�;�ۮ��P�)����h>	%��z�U��3���JM�?��	"��e�c3ކb��o�R!��s����V��D��Ґ�R��Wm}�u�,��ע�p���:9 pֆ��T|Ie	ʕ����E�a�%hc!`7���
�dH���0��A"���� �t�>eDω��Oa�U3��������,11�N�J���q�b0�S8�1J+r�����s�h�e}�>�.�E��gt�؂_������F+0B������o4&��(�+��ڝK�c`M
������:j}���<�ǋq��p�B��~?jv��r�紗������-�������9�x_�j�� �w�Ţ�_�g~3q���6Nuz���J�0���3���=7I���f�j��?i���jNo*��j��Su��ޠrOgz)����v(mF*��(o��z%\�֓&#��Cl�H�#�͉�kGSq �� ����̀^���s̊р�TxOvōi�¶��޲�����U����竑n�L�O��C�<���k@2��Z#1l<��P&����� 8$N�K�_��r<�a���/'�J�T�:&�ˋ8��Z��S=U�V�<daB�ޮHe��W��{G�'{^��6E���A#�1��!6��a����i�����IWm0 ^��s����9Q��8�����e���"�B�1C|�ő��adX�)2��x���D���8:�L$��}7e^�7%�L<z�Qӹ��C��0�i�1��P̛��Eeu�臇�5��=P�r�PH=)�Ӡ+�e&�D�³����,��Q����8���Ϯ$ΨB::nY�ք]V��@�n"	a�,#_3�s�+�%���씦[�W/t������d�;� ��xs�=l����0N�&mN�����-Kp^99I>�c��Y�����%kzc�i������V����^�nr`�ؽ�,
3qbrl1pH�ȅ/��מ,����[���
�<0�o�W"��1�c�d����͞�5d���	?��u�xpӟ���t ~1�X��`ߖ���3ɮC��V�<�Ȳ�,���B�FߜXp�<��yo(<�g0z�	5WuQ-X%%�7͖E��A,	������+�Aη��x&�wG�0-_'��uJ@�h�ҮP��7�ݗ�Eb��L4���^Ѓ��D�R�21H$�C����"t�������gߙGr�����v�G<�|�=�����~�bѺg�y������H� ��-R*j�5SE:&W�)]
 �b[t�b���+�O;�?Sm;�7��9�.v�.��p@,�+5wv{����|�xDGi�V����M�);Ƅ�GJ��h>�h�{��Qk��� W�6�j�Vְ�Lރ%o�p�?�n��qnH��ߋ���|�.L�s��D#U��G&,�*B��D+=*��$��L��?:��FW]�ڤ�� �&a�?O��2��eaI��?C�����z��N~�}�q�AFK;L�	�P��S�g��Z_@9�F�q�_E�;
�leů�C�r\�v�@`��ؙ��.�����T-�u�a4=�k�q~�Z�����m\m7'�Ę���xu.����_ϕ�'i��$t\X��/ʲW�1���X~��H�n�8K���h8�&f�ۘ1����6nD�1�m��zK��0�x7������Ly�o�
�.���]�U�4O��TrR8ALB��Y��'P��@~.��@�!�Jt�n��Mȯ`D�l�S{K�_ώuj�%ԇ�+�Ԩ}�nh0��q��Z�܂�k��TD"��)�Y��K�s�<��&�PM���?�z��ʹ��N�s��G�<��β^Y8h��s�o1�ڮ��=·�n��&���aI�nEp��~��o��]�B�Y�4�pN�0F�#����d� �EԾ���|�� Y>�[�6`�s�����@1TI�����t%(n�j1ɼ����.��#�G�.2���h�y<�L"��$@��ҭ��T.�1�+�pw�Q�d��U���BR_���A!���~v4oMܬ�*��T�.>7J���iӊTrL�i��T�ۂɩ|�!&��T:51���芖a�9�`$��v�����C ���5�o#S����2u �0�' `���K�/�yW`U4�3e\�ZU������K�W`,6��U��!�p�{��{eݰº��v���άe@�׉Y�@�٘���Ӡ&/SM��h��)5e��l�=G9�͋����b�HY]1+�ɶ��-�%
h��0�-	m|>2�.!�Jqw ��>�ڸ��I�ʒ�`s��>����&��������I%��$M<��C�C��QP�Vt����A�(.@w�6+��B� d3��'#r�{�)�z��˵M�r�P��01��6ˢ��MU��� ��t�U:)�O��8��1��z`�Z����<�X�A�|u3�󟎷�%^�6[i�R�}��Tdk�
�g(�?�i
���b��Q��%��W�6�ǐE�bML�k]H�l�0��a!0�Uf,�Z��)#tsw}Mp4�4��Z�d�DM��123��q�*����ۉ�"�?�D}�W�A�4��Q��O�C�b�!4��J�(ze����F�<�R{�CI*_��j��g�rY��ak0�f����q,��(~V�:8!-b�<�@^�F�j&�e!�
^^28��n���+Xy����KRGIq�S��ƚL]/
{bH�;��/Xn>[l�%��=��^]��jl�����|�W��:�' r ���%	s���K��?�I�BW�v@痮˲_�J4��tJg�wV[0����}��f�ؓB遧������3��{Z��w�0�.t*5p��@:�I�	��
�j��ESYa���B��eJ�K)C�͑����vIz�6ƇՈ�èuV�"1e�8ޱ�C|�3��Si
� D�ֵ4��3:T���ߙ��J��~Z �s @d.�>��^MeM�s���oZ��tQ�P�c&��}wL'?��� �i�
��l����r<IV��1��(((�a���d�5ѷF��|��Ó\��pm�����=��q����o�M�	�R9�w`z������g'��E�h�S�2Q<.2�̱<7	
Hf������o3H�nĵ�l��p�K�1��L����p�������nO�).���O�[�|J1,�J���/��������z��+��g�n6�o3QkX����N�nvH�-h�~�/Ϙϊ,CۜY&��r`͈�]g����4�VeŇ��˯���}�Ӥyzb�8HΊ��/�Cn�Ӑ�_H׮�:�.�̼��{���"�֏53�ȧY#TX�e�b^�4|�����ʚ���ߘ�TR�,8�ܥ`7�x����݋nUJ�xVb[NrmN�@�7�=kDP��KN��Ci*Yy���3j1HBp�E��(_�޿�\&9�1#�' ��?U�4�h�IM#��|3>�䚫U��}�0eL��69�8�\+����
�k��¥02�V, ���&T<��������xC5X�Y�)�4m��x������b5GKKtS��B}k!ܝ�"�����^y��R����6~�JU�� �p�nE|���9�p�kJ�b��M���Āq�*�.]�Vn��&tEl-�R>2����B�9`�{�GI����ykl^E3i
s��}���˴.�H6dS��(��Q�q�KA��z�<�b�KOm��'L�9?�36P�|qL�I*prz��Y��B`��g<)�k3�"2�@�&|��Aڽ�:{N/�QP�D��Y]h���w]���j�Ug�+��S�/�D�E>T=�V%g���͌������Qrr����[0у�F��h+�]?
�$7hhԅfxp�����d��O��'�}��5���-s:�C��u����b~�hd7]�bt(���
�<'���w����vy_���/ bj��\l@E�ky�uH��>�������	�V��*�=���W_�H��PA/{��N��zǇک��(�3X[,�_qm �s?c�)ѯ�p��Jq$^��Cޮ.o�t&*�2�&�	���3�=4n�a/Ƅ�M�8�7 ��[��n�M�%�I���K�7c�F�5��H� ¾Ӊ�nƂ\Ĥ�ʭ�X1��~���+��@�{a3X�✧G���<i�&U��M��E��8:�$m��7`u��i�nXY�'쟺�[#x7�῅ �=@&p��|�"�t��]I�&��'�vN�~"�uep����;Y���'H�q 	���g�"��Ё*+j�m���B���Y�����i���HrRc4��OE�I�U=2"����#�� ��x��_9s����6���k:�?`s�'YX�!_9��y�mw	��^%S㒅<G④f���Ϭ�"���2�x��s�"N���Ǩ̩i�W�����Ԯ���'}�q*�|m )MZQ�n����5'��[
1�:�¬i�"U̙n�`<�LT^
�#ecɟ?�z�� '���:q]M����AM�L3��5�g#��:��P�0���e��������	����zV��*�c���+
���7H�*�^-�|jp���Br�2�)���y����I� ]b���L;4�' � �:D�-TU�Z�g�h�����<�U?R�^
�$@����9�dP��_���HߢW�%'5���b�	�sʏ�i8�ӵ�McN����t��D�]oV�~���(��io&��|����2���΢f<����/"�����5C>O�,�m�@�l>�n���l��U?4k���'�������]vk��Q	���f[�H�����hub�#�D8��O
>������H�a���g�����W�p:}� +8�P�,GBb�m��(��5���K:��Zvj��]��19�SFMC�;AX*�X��Ǉ��!95K�h��T�$�_N�d��:�l�N�_����β�]�k|cf������i��I���o�ԛ��x���غ�Y�	�a����9]���@��S�vE��������=��Q|�tװ�U�u�)0�"k������� ��gM�	���YE�4�%�Ѹ��3��/M�!�*���4�a�ÝTM��I�����!�����Q#gR��	�j��VuǊ'E�W�@�F;�3A��{�;�4f�"v������=�������?��{���E�C��̺d~���Sg�ؽ�b����9���*o�.1.��<!	�Y ŉF��i?���0w0�����;�Q�b�	K�60��҃i?��b��6�]�jz"a�n��A	�m��p�z����=����Q�R(מ�?OY,�Bb�`�q�n�I�y�uu��?��.4��D����oS�J0�$�p_~y(+ ��N��6�J�}т���*K���	6��k��!��C�� tԻ�/�Pp�_�j�+�����
�9��������xJ��Q/\�P�H{u�a�h"p��8�S��|��_-6dM9KΉjZ�q���/M�SC�a`����f7���X�T��L�|!��T�����\$��
s=�,k�B>_U����X�<v��ڬWk��k^��dz���Gy����p;n��'[�T<B�k�����&Nf����_KEar`�����-,�v����6�Qg�/sV�04r�r<�����X);*�Y���5��&�T��6+�����l�8ٟ/�4 �1̪W�r�ѻ�t E���J��`�?ϨuP�������D �4!���-�0������ ӊ��R*�o״Gy��3).:�Z5��y��x�̙��,��@�n�w���;_9z�\ꗝ�[�����\w�^�d�m��{��������I(mP���rA�_��-��8���J3d�W$��*N��E)��ON}��a#���w��M���[U�M�����K�q����Vr���ծ�]kb�{F�w�K?���؉��:�L�D�|����I�4b?%��A���7����,B��A����>�y%�����OJ���@�W�^�V�m�+�0���eU�먦({omV~5�nI�@N`��f$ތc	�����h/aX���-�'yB����O�J�v^���@����](<#PPSQ�W�;&;5Tޞ$�l)ä�IE���D��x��̮er��f)@���(}�
ö�z^0�Ej�oL/�-k�b~�S�=C��1[��_��l���l"G�X�C��oqb�srUax_���[[9d<6���g o�Q���{���G#��؛�:��k�D�%���k�N{�E"��{%B�l�9���礪�˚�#�ܦb��RU�&�����X��M	�����*��MAx�������}Ѳ4ځxD�����¼ҩ��,	��޶x�|2�e���f�[�o�
�6%t,���Qg�B/��o/ʻ"�=
�͹�긌�薱2*��)ۚ�5��?���>����];XK6ڏ>���G�[؊�X�QD�XV0���X��,x;ך~5֐���`2*������������yT��B����ʂ�U�����",=���\!��ǐ��S*��Yw�=a`�¿V(j��E��������G��-2�u������B\q:;��_��9�9��yd�韅����z�1pW����*�����w����!�ʑn��FC�YHV� ǅ�s&��~U?�9�
����Ȯ5�~J6$��=�$��>d�6׶�����(Ks�����8O�_�4h�`�c���eB�P���ůÒo
�K.y p�}�v#���h��i䒡�y�����}x����w�~��7��/�ѣZ{�K���q�V�NI�|�Mt��Z���"��b'�J���1-9�FE���_��Q�e�[�� Ńf�l$���B�2~�}��wQ�C�9��?�թ=��P�g:a��A�]�Ry����s�i� Dd�����5Ɉ:�.��Ɲ�{��$T-�o)��1/����1���RFgٹ1�d��� J�lբۀ h�B�ͭ��խ�{�h��(&+���c�a�Z9����椾{��r��"vj�YsF7�c.��'Pfsr=`Œ3�r;���~�N8Α�6���Eu,��w	83�%�$Q��v�*�sV�hG���������Q���G��� �#���ĮVRl�+S~e��!N���l���`����6�6>��񆅮~��Z&�����]�������+�]�O��wR�rF��Q[��-'��ͭ�	�Ot>�D/t~2��
���S#nL4���ü�R;9D���,9�?'#a�ݳ�j���a=t���<���YB�;��) &l��:?�;�'Vw�lї���2�kd�T!�!�|��	�T �F)J�YƎ��K	�B3W�A]��P'+�OJ:�����OX��������-n8($�q����5��\�&�a]�ۆh`��F�)�S�ǩ���ճ�ܱ��e����T(�ͽx (6�H��O��l�㬆e�V��D!{���lpL����\m��D�c�N�x;�D�Ô�"u������)���u{�s�L'��+��	
���F.�z�1�O�����!�Z�Kj�)W.�u��1�+i]�m���<b�B�"�;�hg5Y=��-��m�DLL��)-����Bg`�W"ͻ1}g:g�!3MY���]�H��=쀵r�а8���;ӿ.�?����ȍ8�K�Oмe���Cck�d.[P�6f���*����F
�Ԛ���y��W��Iv#1ʈ�G#3�pD�k�g.��$�e^�XNи�M��4�%��b/����*��U�V��	��P� ]�%��@�6�G�զ|^��\�Qw��[P=��,I(�!�KG�]c3F�lvR�1���^���.� ��K\��'N�F8k8�O
�:خ:���[aLW�4�~ּ��x5!P6�^�5��ވx'�ѥ��g��rՉ��O#���x J��zy��V&�B	`$�1��_��<o�[5X.����xL�	F� X����/��l-���&�3*ǟ�.Yˠ���2w6�E��l_Y�$-���`�B�2r�߂��Z��/�ǌ	TB�Aܧ�X+�˼V&�WKUF~[c�B��(���EG��i�@�e����wmk��ѷ�q���)y?`��; &�	K�,MQ˅<\�戠}9�>�6����&���g�i��C9���d�Tq[l/a�~��bhO�kI�e�O�����9MD��v��&���)��SD��!k�]�l:H��36;7��,�dm�Ⱥ�K�Whmz�lC�2�DC���}�Y��ɘ7_g��#8H��u/�"[��`���n�>�����K+��M��Tp���#����)��2����Svc�+��P��m�C��֮8DE���V��<.[��C�E�1�%s兇'�㰻�o� Zhnm�2d���EJ����o�T���کP�����S�ӿ�����Q�˹q�7"���|F�F�>;5��.ٚy�F��'ݒ\K��b��y�4C�L`@M!��G�(�Zbr?2�d��aa^ �
�P��Q ��,$>m�P��f����纒�T;��?s��"��E\.J��K�]��ݣY�����ɠt�$�����d�|Ƨ����K}<+��$%��UXa��ɔ�~c�UK��/ �X���n��Y�-���I5R�z�m��Z-�
�X/R`��6�~?��X�~[����LJǆ7�,���p�8��l:)u:+��
����tk��4n��N�MN�֓&ͧ��'y�_�<�5B�Y�wF��1o���wt��0u�f���$7�L���ؕz�K�g�o��������^c�1��v@4���[�{S4����C24������(�v��/�;���xeW������t�av(�c�?%nm_ �ֱ�ӯd�(��4�C�L�y6;B29���,@�� z�&nNŝ�TIh��U]AU�!�ifRyiH@�:Lh�v�f{p�R�ҝ1.q/{l��a52I�	|M�_��
�0ڲ����"A��Y�ڋp��p_)L�ϑBЃ\���m�J�����N�O�	u&
��	�L����K��8"��n��-���j�{��k�L���{@O�Ef�Ӂ�C�B�tB����9sV×��Ӆ�@�����L���[����O{��ݐ�k��]��bغϟ!D,�N�X�auw����+������=��9}�\L4s�}۳��9�H}��zZ%X-*�!~'dT�i�˭JK�N��j�<�b��=�h�YL�t��h�3ҫ��%Sp��p�}FK*1I�.P��*��r\�A��Uq��j���0}��T�\�MlOh��t9�$����z�r��%�:"��?�_�b�k
��Q��}��n����ܴ�TСU�

	cg��X@�h'o1q�����0Mc�$o�hW�N�L�6�h�*|�R�L��NY�ă��|�@��p���jo�G�}�#^C5�51��r�Rr\�o�]�6�c<�sY�ifj�ӓ�Q`����I�S�a��?n�\5\� FZ�
s�	3O���[[�5(�$;Ľ�@��� �Q��˥R|�6@���7㋄B:��	�sD0Nnb��ʾ��BRh���ZJ�9���Ԁ��w�U&���J��nԞ��T��
�I������v���:�J�nW)�P'��t
�+x�r�2K�t�C�}2�mj2~�����/�!�,���y�d��|;���[��>�fJ�^$�i1��`������+1^|���Lbh�za�����H	�~��S(�}ѧ�\���Յꨦ�FD����L����%�Gdv@��ҔY
��]
��䝒����<kÐd�Tp��o�H:�C	�-N "Q�t:�c�2?'(� �~J��F6��C4;/i��Q���5�Ȏ��G� �ԧ�Ȥ	]p_Z�h���N]���_�B�m*��E��Eq�:a�;"(�6�a�&_/h�A�j�ApssV礪�ⳝ;=��̓����2�^B��!�}�$�*|VQ��:����06��>C�]��n�wO�]���TbV���}Rp�k�橠�즹��{����z��]t�^���/���D9�fRSF�����z�_x3l�~".���\,E���)sz/j�ZF�_�$��}c���|F�t0��
����'�A���P��hy�G��	J\��T/�W����`������j=5�w���^�Ɠ^��""����HْE�a�q�	�����~�vTcK_W4kp~{d�tB'�����{I�\aq���{��И�_�D������������a�x1��OZ��=<:O�PZ"����̀���bl:�;�^0{7��sK��J,r�� zV��]��$q,t f7�ҹ����稴tOa��������<��+�B�j%@���i\����{�Pm ��e�0��+��i��;��Q�I�Ee�5��=����:���=2�����ù���_5l�_5�~y�{��#l�=��Љ+�ǁ����(nьؼђ���w%��u[t�Խw�W��T!@�%�ߊ��8CJ��WN
�I���t�^EO蕨f�X]Щ�>��.�EZB�'���4�T�/ޮ�f�.=� �ބ���;!����& ���؎膓��� ���(z��iDŰ�����dCe��w�Yҟ�[`�r��l&��-�����e��p!`�ξ�q���+�q9rU�l����d��bXL1�������4Sƥ�&�ʱ�h��CoS?6X����C���Q���-I���ߞ�wh၁��݇=}gO;3L�H6�3�E�~���f�O|���68M�&�çEu<O��8-��D~n���f���7���
g���QLu��,ġ���!f�JJ������l�%�\Ɋ�[|��ekw��;@�n-��H�x^��	��$�fR�G͡>�-t��O�i���t(��`ZJ�F�/��V��X
��� D&xA�̪+��o�Ƅ�GlQs�`�V@�ۨnĄ$>��""�I3m�����uX�p1�׉�K�o�Y�m�-0A��MN�Mg��#�5�*?���{aq��q�9���.6M������!�� 0�㽃	���9��&`tO����{��3ʏ�.�.�R�F������r�sE���y����ÄZ���P5�킜�F���JIv����~c�w�>���bue	�X�0���A=��y����j�y9��O�w;�Ӣ	ij�+ �Z����u�}c��c��@|E�3��26�X�U�A%B��nAX7�[$�E6G
�q���޼E���v���܈�k�<��X�~�-YUG�`&	����ض$�U��bA�P����5�G��C�Ԑ����K�8u��fA<}�O�ҵ>t�}r�~66NxSD�O����f���μ@l���x�3p�iPꋳ��
$pe������*��M�l���$KVq#c��;���1��[��x�c�k�P���cb�,���<3��(fs��\�h(��Z{��nL�FO��K���¥b�|ޢF���˙���UtB;���{ܷ�q��xhnɋ�Vb�x��C�l�EjgV�/!�Ӣ��0Y���E���Z#��Z��Ŗ�wĩ��t�G��|\�S�i�v $��T�V�`�����0����/��{�I�glGA�Hab\'�η`+
��]��.-Pq�$�4��D�c>y���� �(dϠ�g �#b.-O�alO3���շ@��df�?~�A�v�\b�gQ7�f�r7��Ћ����Y��w-�j�aЍ]W=��'p�3���O�����Db�v.-F���q����hm�dA��p����:�7��t�.X��7L�!~u�#;���$��ԇ;�o�qzH��*m��ԫ׊��*|;���!���������p��⽧Qm8��t�v�*qp`!��Waj�r���6F�:UY+�t��q�h�xyt�����:]�4j�R*(P�+��0pHɓ=0)��XC-�R����� k޻q��M�{ZL�*�p'j۠l)���j�WB�JMف�7)9��؝&������T�.���嘈��/7Eǜ9�T��ׁc���o�z�ծ��ӕ�Z+9���}4O����>9��Dt���E`��jz�� 4�	�E�Jhl/�л&�p����kR������������!������1A✚da&�0�Bʘ�� ����y$��T��ɦP���g�gr[�H�p:��G�rN�7��^@W��6\s�k���8:���Gd�ʷ�3�/���j�/-w7���&�o����`���exv�dP{��c/Ci���(�7h�i��l^�8��`�uM(-W�s����Tp[�Ď�K�R�`�F��[����=1j���dܟmlL�_�=��xzf0��0�O+/�tD��\
]O��_|�j��$��*�7�^��rӆB�=/F^0��˝��
����+��T�/���ii� ��8Ԛ�^
�"HC�>w0�rO�r��T?�� ڄɱ�&~ka���,]��h��ha��S�����0�>��ɑ��k@6��kp��_�YĨ:�ϓ9�u�CK�<8,���$� H���RDrR"F��g��[��Q�T�W�(<6��
(�������FEbjwH�sn�>b�����fs��:�r���F́6�!f��������j�O�|�3��29y��@�sAؼ�S>�C��pp�Q�?����Px�/��̄۫�1����O������\�Ϯ7VXI)&A�VT�<��
��u5I�o|2]�cK�(`�1���3B.�7��Uh�w�oHq&�i�zvm�T���)�t'YuK�B'��H�eN�0�C��Ѽ��@�О�,��Gn �>6��l�"�RH��k�EEL�D� ����r�!ź!���(���)�����,���P���|��E����Ya���[��dƳj����AUG��k���,r��t�nn���l�j�K�q]��7�y;���Ni�����Q�#ҷk�Y.�!dt��D<&#��m4��y���;��쒧�yY�T�7��z�8�&�Z�M�F̫�O�����L'17��s��aK�J���nrdB��u�j��zE�B�ʦ�0���m�wx��?�Y`���=����]��gc'�<~�wz$$�����qH�r1UP���-R�_�*X�\���ϡ�P�P�k��y]�`Ŷ/���M��V�����%/>��ï�V2����rn����wʌ����o����;]>/��ҽ� �&���,-���0�z�����{?c����>��Vd�A��cɘ�ߚ�RϿ)V�1���w�<V�쏉jdM�e��'�`�>/�SʜI�)�]"�0p���ÀXI*��'��Sf&-���ڍ��F�Vkf�Dqo�z��*���e�)8]�]����1�p�:��xV����Vwv��R���6��sd��J4�$�P�I!�7R�A//�(�(�GPi���dњ�]6�cT���8#�-)�8�����X��sf������92�O'o����iÈ@�n��
��?���hl���u����t��zg�f�UQI��R�;3j��E��;�������ƀ*8�8�/���k:"{�}�+;�E�G�'X���#<S��q��'�B�a9O��W.=����~y�r���r��~��򪉵+$��!'�����~S�(Md���u�8����.�8�
�M��T/�p�l	 ¿<��?�A��?{Z!gK�7����-��U-�\=�`;o���0S�?D��:�q��y놸(�&H[#�Ym'�"m�3�[��\Z�x�u'���������uޤAZ0�Å0�K&����� � ��E�l�j]�a�R��"2�]̦�B2j(�&e3qJ�h��4�BWq~�c�%!��6<��MCd�A�u�Y��+�2Tj�2�{r�w*�N���x��߇���gy����EY��F�Y�����ۢ%�Fé=���)`^q�l�k�yt���LɟY��Noؐ��d}�*�P�03�3%��o�"������$�A�`�DW�V2�(ր�E�u��4˴�)(S�4i0������/�3�L�@#%�C(��6�1
���W�|6ٸ�VE7���~��[�t��O����a���%R�-�v�0�%d��&S�5���wF�x�-/���y���Q�i�CB����Bq�����]�Ji����"�A�B4�XW�������~�I�)6��|� ���u䊠�f����Xԃ���K�*�n�ޟ6��Cz��v�@
�
{>(zuA.|�d� nf���%��C+�mp��o�)�������D������늩����X���[r�K��|||4y�*�c��<���O�_�����f�u,����RB�x��$��M�&�\��}�z�B\�ː��d�����|�Ḿ�q�wAؗ-��=�"�:;�+��'M�7�i�;��{$c�V�M��������c���[.m��o�i�#�U�������PV�l�e�����i^`b��r$�����t�Se~%���(��@�O@�� �d �*2Ka�z�,��2V�"����a��(�� �Jn��� �7�T���鄌�m3�>��j�5jA�IH�6P�B��kL�;k?%�$h2eJ��Ł���W�1�{��ޜ���\�b�lh��q�5u����$y(_�ӿm$�̖��X��¼	Y|oA�гi�+�2u��m�H�C�[�|ܬ�Lڠqퟞ�޲���Oi!��7�|�{���3��Y�k6���E�ILp�Ik".��]���iO�ʭa�S��A�Ta'0ǰ	0����eY�n�Tzs�%3��
0��'1������3y�`iGO"��"��GY����r��f�>`4/�����U��D��yK"����'��l"�\����b��A��WkE�<��KOM��6�n�F�x����z���8Kd���5C�w߈2�xPо���n	d��Ff&ol;��>/�$t7q�&q���H��L�hP��XvTRq��	{��@LE@h*���f�Z��'�<����dϖ�>���E�m|
��+��lJ�T����)�Z���P�/�L��\�N���c*�1�0@|��$w�9��M�1��&�2N��+PN�������hyb3�G��V�T�_~��X�؉���㰕	�9����-���NGF���a J�Q�r�hqP?q�!��	7�؀�DL�Ú��$i�Ɨs���o�&���f��kO�U|'��\C�]^2!{5'{��Ss��dx�L4������&��n�/�a���=B�����#���e*k"
�v��R�X�5��~Q~a�nm�r��8K|I���򿍎�����psa[���g�-�3ZCZ�<Pq�4aH�5��A�F��U�}YsR��CE�%5
lI�(L�F{t�KA+H|����0�b�m-M۸�W֒?�dLщ��+y�R
bc�' }���6��iı��-:ʔ�4��-���<d]G���s�|�ԓ��ȑ����F9��J��}@��n�!0І0�X���䷐e~}�V�T��Q��9��> v������%ϊ�6m�`����^"�0��<�K���@hkF�3����jsSj|����V�w�I�	e�T�Ƴo�N~��{ԓ7�������2�j�<�����.l�/�5Y+=7�f�<�0LGQ/>F�����p�4��	}HÏ�iX�M ?�q;����
s�Z�j)<��^I:H=�"ێ;��V+�-
 @�VlZ)�} �a�7�(��I'�;X�/�N����F7Fo��(9����bP�y%u_CJj�:+�2�uc���s$�I=s@e��9�;���[ٌ]V��{���H�����ͯݢ�%��T>+�Kb#��w�x��X!��lD,�KX�6lz0�z<%.�o頩����REJ�	u�乘�@Q���L�o8��XȾ7Z�ly�V�WzO'X���"L���[$;a�Uܡ��w�G�4�BO5ۘ�����\��pIha̜��-�a��3���`03͡3go��¹: �b̻������1L���v�,kU��GX=5���G%��M�X�F�XRd��s��0�H�Tg)1ґ�ga�lFB��k��w����<#q50e�f0u3V������=�*+�?L�!yU��F�W��r h��[Z�,(3v�:IJ��s(���(��Lpͣ�P�\k�]~���F�V` V��QNM�c��˴XE������{�v�[ӧa[*����:�@�����'c`r�-��� s����I]*�'�l�`Ċ8�6O����#Z�tMn�rb�b.Dw��k�Q����<Z�^����|"�׻p�`.J4�ρG`�����&u�%���+������t	o\IC�����n�F0�E����%7��hZ��*8*�	,��E�J�8�Wf<9�f�S�ބ��d"UԤr��]V�^�5c�9���_Y��P�C�����#r���=��nelR- u�נ��]�����gʽE�tY�t�J�[%?�{�+�������;}Ts4:D�����$��X�C;��=��}��b�ZZ�pE�y�0uo��aS�z�M�D����/<a}�Z��]�6L��.�M>��n�P������8��Vq�R�P�`����2�n���մ,���5N=����d@
nbB�ۂr0*�_fI�T�3;���Y׉q�2�u;0-9k�B���x�T-��Bw~J��z���5��zU/�FHG���	r/Hr��2��(	_���}��q5�u���kŨ�|�V[�@��}SJ���%�³Q �Z�6��`�<j�.wk���4O�\���&���?�F�Un��9vT�Ys�j���u����Ca(� �8�������ISk�K�Ϳ��?��4��F.��|P��� �B �Ӹ��J���V��7�)/Ee�ɋ�, ����|s�-j��%��k-�<ܞ(�6�n?V����c� W�4Y־+T'��j0��W7![Ĭ�#p\HѶ숒�.���Ф	�i��b�cݿ؃���fP
��AO�T�¸T���h�6ct��P}�������f��`ޅ'H�L�U4�;�(���!�]����xz��kc:
���V�$�@�X��$J	��FBE�&�`_}~u��f8Е�Fr���C��֔H�g7�,� U�����G�i��V��%%��Y��ȓ�����?���V�.�>HˊG�G��8{��ڗ�'�?�M|o�r)Ⱦ�T����R�M��Lvp����b���|�����Wc��6q6��I;կIbh\͔�g��.-Ƹ��B�i����� ֺfgA�ּ�ZSh֦q�����/n[Z�?ޚ ���I(�C42��O�P�#�����T�~�F<@k<x;O_%�y�ݣu$�'�[���kX� c7�UTFk��9,V:�CפFl�5Ymi�	�&W v���hp�5 ��A�"�[ԯ�5V���q҆�/����Z��v�\�������>�U�\-�<��55��]�.�#U�,�I��:meM,:���mZ}	K3�|��y��6��lK��������+8m�h?��4�O��w�8�����Vs-!�x����^�Vɍ�[蒙I%���lN�{�g�J�J�_|���-5>�O��ش7�9��0,A�T�������Hf\�ݾ�8!�a(/���/'Q���x�=WA�5 ����'}��N�V�q���e>-0O��_Q�\k�7�*����l��̹? �� *P�����H��e�ȉ���=���8�o�(c^�l�YWh5��)���#�����jhiYǵ=�ĖK�\��L��s�)U�!4Y��0/�t3��b('-A���/_[��Ӝ��^�׻k�d�Qm!��b/ZC�t��OF��	a	�X�hǝ���&�T*aWt�-.�,���L�۝:�i^Cn����l&�b�\EI�l�}�)�e� oN{:�pO���͉�&�β:��M �1[
M�{*=�T`�������dw��i�D��,�w��#�����l�x�tz���&���j��6���6�n+� �B)0o��5�@�e�N??1^��Ｙ,&�sryK�f�q��9qjCӝ/-L�v�0��7vw]܋o�� I�eP=
�s6��wni���}�v�4���S�1On5�O��X���~���p5	m~�05��Q�0�Ԉ�-j���%���߯�`Q�uq_��bF��O����R �3�x���I.����i1�\���9��Ut��yDJ+HzF�5ݣ[.K�Ԡo�[�����|;5�Gj:"���Wm�w�sc��Ȭ�5�"�[�}T���z0�*�"hx�����1��y����[��}�NIކ�i57��N��{E�庵���_ײI_��k�����D�NP�}��R̥����p�d������*B���m0��[p�+�	����9Y��(�b��P.sw�7"`���~��F�2׃L+�K�}d��_�Q�iV	�q�>ɜթ|�]���jb�˱'�a�I��m� 9�gm�t�7�^O����0�����b�P���=�'G�ڶճ���i�~�K�M ���_��=���$��§�cO���i���d�mۆ�T��w�Xu���sa��)eXqD��o�ڳ�]g=���Sc"²Nb�8�Z6��>S4��xRP9�tq���nM��2Ês��7��B�5fyB/�\�K�aK�F�.�~�Ŭ&>]f�І������/y0A���$�I���.�6��u�1�VN�4~c�Z��z�&MB��[Z�a7��~q��)�Vͣ�}�l��(�0�4��C����͊Arc�/d?���&�ǻ�����Ŵ����|�r$�s�!]���?�������.Xa�E3/1.,&Y�4B�y l����Fz�����=�M�"�I<�N��𐈍�ٶpu�6z�����J�y<�1��L�A��5��Yc�[��KQ�����x?��Bqu~���y�`ŵ�r�=a�<���E�3(�J��7F?�/�̪�*�DoTwn�J�$�u7Vï��Mhp?ҟF�.d)���o��G�?���a��%j֠ː�z�@�?�P�Q��2.�	)eNpű��˳OT���n������SED���!�x�UȒ�4:m��Lf�v��P�7��e39�����4~"U-0_���0N1"Z1�[������%o�'eN �Z�z�! �x��-0�:��ek�!��h����[�AȞ
g�[jp��r�c�K��{ĠƦ7���U�tü�̓��K=u	+I[8 ���\�W�`0�L�����d�yc̏��s껎ac�4n���J*�e�l�FĘI�1A�żzQ�>�o�Ǡx��H�O���ŉ�tx��"�t��1�uƲ&��A����*1�
5#�y��6��ZSX�	x��"w�ëX�U%x���ˏ�B�&-T�
x7�+�֜�ބ٭�(��I�pIj1�)#h�O�G��=!$2��1�8�i L�BH8u$�=f,�`��z� �%�F͠:S��E;�t��@`D.��(�V���Z��=^^/A�N���M-���C0����v�q2	b��;jF{��}�%��Q�$��x��!E�'��Ү��_ �32�]���@��<�3��	���M��s1A�ZZh黎�#���*lٛ���-^�5��Y�g��Kᰚ���U������?<��]b&�gfW���=R$V�Н=pt=�V5�ū�0��	H�<�ūuY�U
àz��c��e����v�Z���ш�B+���3�G��5�K�X��E�9w��@��.�����b�m8��}O�y��T��O1��pD�M����N<�`87���봹���X]&�$n�Wu&���4��,!S"}3�f��<�72�� cߊ�òr{�>����	Ё �@�Z��ԁ��݉a`�`�5&�Ib�6z wb���xsK��͍�=
��cpӉ�pˍ6�����q��zdh|g���\0>]w�5�HU�7�S�^�CgMA!�Z�gb���5���^C��
-�}�-o��I�������[.7�Z|���e�| m>�	r�46>p^AP����@�=j睹B���z��Yic���bfV��!Z�x�Q&�}����q.t�Q���?lX[�xr5�Վ�0d~����ꥪ�_s��r��Io`s=�3�8���WɝT�nK  �����3�8��i��QM<����k��KKN�HM"a�ӉY'6~��{�Wb�l�P���x/^_�f�u?hP��_j�*�2��g��}���Vaew�WE�=�y�8ھEH�AX7�zv.�J]����
�L<�Μc�hl��u<ԛBb��;�����^tRm�g��WdgǆF.�uV��I��']�m�( X�+��g;ў!�4M�F!6i�FV��P��RQ�}�ç��I9lL� �Տ����]�(͍� �dU�5��\Un c���?� &9``楖`�޶8ޒ������@5�-�'��z�yZ��	A-KPF�E0q'�����Q��ęK�/|B���Ldl��R������i�Go�o�=Wy��	���,5
u����B)jì����/�　sh�V�Fi�*��:(���5:����^�2��EPd-��愃(˾nQg��4��N�;.��>vJ�O�� ��az�J���%Y�T�CS^C�9����Y���gR���6�Ξs�~�Pm9l���Q��T��isu���e��Y� �j�_3*~����?F7�;�f�i?}5��Ǽ's)����mq��O�JݢLMK�A�u��r`{�~�[mw#�;�\�'}���e2 �A�򏵓M���7½N���I��a����gc$��9y��i��QY�prO�a_(h����&Gh�݋���Ubz�����r��������(Z�Ԝ�=�<��:��o荪�3}G�����W���D��WFؕ�Ԣ�7p�u��a�Q��S�\�����~�#&��f
���H��ث|�C�"��Is>2��K�o�*NY�7���ܖ&��#�|숒����L��@�ʸ�X����m�w��*�\�1���)u�����g���ew�8�&��Ӆm�c����i~#�
���5������u�2�����V�fY�e��l����ѩ��E�^�Ľ�O{���c�CZExK?j�}���=�="E2�.�W~K�N�J�G�:	SߛCi"�̈J�F�f�� ���6��
-����Ͽ-^�����݂A�����2M�0��~U^�9��0����eGq0���Tt'��P��Ʊg5Z��u��1��+��!��`�H`5^�[y���(oV��f�p(�ѫ]�,�bD�<!�M:�O��IF]�!1�(Bc��BT|�5�����sy�w���х�3�nIUtv�:��W�t��gO�֝�0@�|e��[����ƿ#T>��]�`�!�k!#ǧ���e3�uU�}���/�L�fu��Ҏ��%Q�	��]k,;\.��Sn� 5���kaD*Sl�R��ޠ��e��yAUb�މ�+t�c��� �iD�n���S2	���@�"��08�y�/��*z�F��L�D�G�}�1ݓ���krA�R�a�4�֭��'�"P�/��M����������C�.S�F������0E�'��`��Q��V����1������o0:ia��y}hp��~yŶ�N"R��އ_�3�o+������V`�ј$Μ95��f�u���k�yp�R�d'��d�1_jK�n��rQ|��(��w���ʰM��_��|�ʋ���'i3�#/V����d.��C�U�� 9�jb��]�"A��N2�ˎ�t��*t��Q.lR}�j���螦Am�z�8d������Pa�A`o<
�M��T<	�T�>��uB�<#Ϧ<K�|Lሳ�'`*$��a��D�_���.��h��
����L�-6�ڂw��qex6.&,�[l���Ҽ2]�����B��0�����+��!a���aÔLusI6�-��%���1�tI?B3Z�����^�s*���a��a�"B�7B7]����G��(�~�z���T����#����a�{����X��b�,?0]�� ��lS��'�������	�WE(j�ZU)��q��ş*[�:�_=���kU��w�K��p�{��b�?��ϲ @gVu jA��]A���,��q����i܃K:�����ii�,�b��^p��K��
]Ibk�zé��L� G�W��q1	�\2�����D��4]0�G'u�ʀé����WV�4��`5���"�TNI����Z�o��M�j�Y�����b����U�[WGK�y�0�so��ׄ14l��^�_�)��W��V!�:N{V��M�����K�4����kp��������R~��9n`�BO	�!d�����)�.���h��	"!��|Z6��jo/X��w�����O{p"%�d�I[d��i+}V�00,oX˲�#tAв�]D���%��Ap�܈��Fm����#dLM�
q7��w���E5�����C��#�tl�a�x�r��റ>�L����ӌ y����R�!n�����A��-x��X�u�2cg\���I"�H=���n!�b�k���k����R�KIe�3vɵ2 -�k�#iS�(���\V�%�FD��+��s>򁹻@73�'�*mH����FP�i�M{���ަ5����p��J6v��Wm��g�b$�/�v�翲
�}"��ɳ���Ai�ݭ���B |Fgk��A[R}U�����Y�U�4yN���L&3�����ȥ�ԫ4�%lY���g1jXT���%��)�/w�7D��ɠ�cX�W<QoA�h���Z�x\�ӂ?ꩇq��?�eӬ����ne��g�a�H�tA�����ዣk=D��k���st+ջP������PZ!�A����'�s�T�8��4I=
'SF�ˠ��T�h���U��j�af�f��s�4���y� /�u����`�{Re�4��w)�8��	�1l+�c��ҭ�[~�-o|O�nQ�=<'��  �r�ͅ�;4d!�R����}s��]���m�em��f�{�@DN�����U��D;�W���bK����avP7�)lv}�V�_M����-�C�ߥ�{���9ZZ3�M6ߠ!� �ɇ�T��U���2�R�h?�B�? �G׬Y_|�]-�6��ey�٢e��-��$Ye��(͊UB�$[�8�f��t�r�!{I�_J�/7.:bq?Y��sSwL&�&7D�.f��:�8�K��ۥ��4R��]`�5/[�L�v�6��k<I(��
���g���;�y����i�8׹�e�����ҧ��p�ԧ"uyk<H��$W�m��-��'��]�f���g	%ח0ƀ�.j���D�w0����!'% ��QR�g;g��i�<�u�Qx������qv.�A��/Z�� $N����I�uLO�q:�����s�@v-�t�z�x�d�o�+���.�=��k������j?6��g�����h��	cWw'�{�iQ�X����$g�k�)�.%}.��"�qm��Ä�ܢ[��;o΄	h��gF��N��qy+�N{������I�1ж^2Qh�i�]���M4�{iۗ��N�14�k+GP���+s}"o�G W�p���Vܞ�2����}y.J�&��#]9��I�PJQ��ʒ=G�Y�[�U�u�s;�)Ҍ^����/(a����QuA4�Uv'������{}Z��3���l8#�ŋ�l��g�j6�\J�������=�h�T��o�c�`�#����8NÎ�M���}\��bb.��6'Hf!&��ͥ������Q��dRɽ��kq�ԎOe�(A~���+2ié<���6���|i�����TH��,�ׯ���(�d;3>�k3XyU׽j���M*<��H���O�d�[3Ռ�a���E�3�"�i�n�~��O���B0�����~�`����V��h�^�1n���MckW�
�7v1'P5�� �a���3w���ܽL�(ݙ
�~�\��{}E�=�r�u�'5�y���H/&fN���݋΅Gz�v1Z��@#������`�.�E=�d%V1.|<�'� U�婺`��$y0aԢc��[`��
��#��Y����岢k]E����Fg40���!6��;�ՒC�g+���60�u�|ktrf��a<*��B,=5i���t���,�v�;�4Lt+>�{�����W��+b��edW|������6�8�Eg{s�����Eq�0pj�_���P�)@�������0��b��P�xJ���+� ԅ���^����Bb��7*����1K,E�Y>u�<f���25�$i��e7��c4��q�<b�(�V�m�V"=��d>s�=4	������P��k�"��3�W�t�q��sl�^\m�rh��3�Ԋu�|2&~�d$ہ��$��DD�4�UY]��F"v8�9���/sgY���޸���h�>��"���lcF����ݹqf�`�ʹd�&�z1��y�N�S��T�\x�``P �EJ:hǓ�ߠ�=�V��Bn���J�G��֣fJ��}� �K��!��$��殺ڂ,C�
�<�2#�9n���S�f6z@z�5��g+*vݪ���>�y/�{m
�u�Ω�V5����߽s�����.U�P������(h��Q���$���\�us��,У���Sq��TY�x�)J�s)
�&V�)Oar^E,M�wP�ά���(�<K_q����H�_�D��'T8�"^�}gxN�T�)������-M�]�ř�ˈ5a>�s:� FNV�%
�P��8��nhq�A��m�HH�Z����$":��T�b��í0Ӫo�X2%�:ػ���"�O���_�k�O����^��1YU�޹gqm2��x�+�ꆅ.��� AL�ڬ�vZg���jWX@d��lu<+hԓ��s���C�NPe�'SVY�昇�G�#��d���6d�S�L�D�#9�q������j/G�b�5�bW9�I"GV10#��.�Y׵t�x6}���#a	�<�O�⬛uS�k��u�s3&|�'��^��p�PH�_\���Q킮zx,�������j8�,w��t�e7	��4>��3�N�ޝe�j�+��ɏ�Eb��b�zq�y�py�x�n��'��/�� 0o[G2�/1f�&������kzf�u+W\]���Lb�yk��M�����a�n�2t�ˌ���u��^ �֨�"b�c��=�f�bX�'�\�*!{�]���594�|���x�/�o���ZVV�/�D�a�ϣB�S�*����:�YC	K�趯uSB�3�����
��S�{�P˗�}�,{#��F�	��	*2��D G�Zr�3��)���� �/���2�YF�3,�,y�A�9�D���`��3e���ܔ,&�`g���b�f>��8aG���n�K��(܏��.T�i�ɖ�~a��K��]eN0Ht2���"`vK����3#еu@v#�k"�/�B5����J;v~�_������u#�9�V`	���L���Q9�8�d`��8�7.���nY���݌��}�l_�<�#Ա?�$
��c)�/��	�� ؀�J�!�t��p��&��E�jJ�C�R�����&�%*��ܮ�����@6����j��{����N��j����#�_P�yK��5��
���D�r��u�M���q&ʔ�/þ�0�o�t�����/+��8�V>mjȹ�	2���q-������j�.�T??F�|N�J�aP�`���]eq�Z��'�G�
Y��.�Gٺ,k:2��_��ޓ�����̅���z�z�b��y�+�n�V���j��`A<��s���/X���>���Hֽ���+�-l4��/
�:j0�!^�obIi��~�gB�n�=���77j����D�̷�Sz������1@iW�!���Cs̾�)SD�[�1\��ځ:���	������0��M�_RF��|�~�-�9^7���T�)Λ3�j��+����ch�*;וּf�~���o;94R �IN_q�Ɗ�+L�9�5E����� ��Z$�9(�c��$`��9-��^żGH�ju8M�no�ꛓ����05�c$ݳ��O��a�m�6��?��hk��\mI��L�(�߱\L׆G�vP:ǘ+���i�O/s'nn�����܂G!YlD]�W?m�X3��b*�x���?H��k�$\׾9.לE�+JA7Q�|0�g�gt���C�τt"onD��ִ�������Ll���-=�Ԙ�U��`��1����ѯ>\W����}+�B%���c?a��4����Fǵ�(�.�'"�M3���;�����䞁�2�Z�<+Q*�w�����(X�m�޳/y��?��uP't|\	E/!L|ܔ��ж�X��Ԟ8}7B�Iq�T��`)�x�U�}s<";!T���oC7������LG�Δա],R�RN:�qCh~X����ѷvF�1-��#�#�z�9I��ue�i��y��!����u�<ː�(�P��w2p�+��T� &���D�T6���c��Ȓ�-\�w���^��J"�`�)���3"�A�~ż�����y��q������������
P�X�g�&ǡiH��}tXI�Y��ǝԆ1��<>����д�2��V�i&�*�|jb#9a�{�����
#nqw�M��?�`15�v��W�Q�Z[�_N�\n���C
��t��qk1�����y���X�6�|��ͩ�b�ke_�u ���`!�v�	恢ӸrT⑸��u$��?�[U��A�31����8�o�w�B��U��Q�ꫵ<9	�ʚ�H�3Rg�c{Q����j6��1��N��Z0r7���߬��0�\�����z�d�cA&}�L)�*aEX���+�]����t)���H=M���v���`�-k��;�!���i]6	
��]���|M�����\�����}����޽�D�ͱU���q�P(�7\��pi搨�g��\k�Ew�:f�"�7�2-9#"'$��Ay4��	���A���˅ZY�A�x�����+!bb/��#<�h��`b�L�6��x,�-����HM�U�)�A�4�I	���ƿ8#9��d�p�}5Ͷ��j]��|��U�ϨV�.0�׽���������3[U�±g���'�ɄK�n���/9�(�<�]گ�}�`��nܯG�=����wLy�w�-�~:d�DW�Ɍ)Y�l�<���ɱ�
� �
�1���W�@���D��<���;G�d(H�Zy���".�aLV�Mf�x>Wד�pJr�{֊���xJ���Lpqɖ�R|�5�����&��k�VT��}w�S)p��:�v��~�*~`��S��*�}�6#�����ȸю4#�U�'��/�[�����I|ݩw���Hr��mˏ�A�d��q�d����u����5���z0)k�+xT=Ub����_�a�ǭ&�y~���hN%�
�Q���QD�D9��t]ĵ����������� �3�	6��^5[+�����;t�V:�ն����W��%&٭�-w�ëM;o��Q�T�r�G��B�y�C=�-�1��%� d��,�N�r�ֲX�9>:&��/� C���9E���b������Xio�+�o�\��+
%�vu~�:V��9�����BI�H��rʌ�K�k�
����u�Ħ	�jB�As��B���H��" ?�i�TD�3�j��<?�lzc�@K��n��Y�����%N_L��S�nu��Q�����>�!���A�H6�'ZG��4+t�2X�{$n��ym��]��p�5>���y��$�+���T�O�&Npp�'_��"�w����+Ǔ>��{�&p��cO�r��}�T��0��&�a���R<e ���;�)eܡ��t�.� �Yf6}���{�uP�m������\���Yz��h��<�	Ծ޵��S,�x`�����p�\~�o��z�i�p&{�o�It��2N$�c6�08tn��`P�Z٘t��1�?����	��J�����]^y��z��%*U&T�����qN;�aH8�6x�W�9����QUQ��>0�#̰Rګ�Ը��c;9:]n��4K='y�H��S9�#�F�������?�P���i�">q��t]�������ݨ*ъ>i��r1�TH!����N�[�(�����30��t��H}���-��5�ml�)Z?Wi���+��z驭QXS�?���ڕ����-�,=��g�G�����%�/���N�4!}h8;�Ǹ�n�haQ�f"S�+�w\�����B�m'��#kv�G�Yq�G��Q���&� kB�B�ED�h�A�����¼�����\�I�w�q��M�,�R%�%1������kZ��6��7�t�4�8[N�r+�ᝦ��x�k��9�܋^��Q8 �g_�Jfu�E�dl�f19<j�q���
T�A�ƀ�:��&�����" ���0��s*�{��b�N@�q��oTWR
�4gLR�Bdk�eB��{xu����s��� &�i�>9a/��@�=[�����Yl����3M\����n�U�!�o�����36c�����?HJ,X9N������>@T#|��T��8��\����aEd��v�hR��X�I��?d��T0�ַE�mDϫYV�9�V�]���ⷡ���g�q��c	�KM�.�����{C*e��ș���w�J��W�7w�x�	}$8zF�w�B����\<[ �0W���2*�&��x����M���&L�����I#^���NB��Cp��]f	��0��\��V�X(��/Sk�@�?`T�0��m�@��B��[���u�����	�_6JZ��8�0.��t%�ƶY3����M��,�N�P��YyJ�Y�td �.�cˮl�2���9i�O)����;������A�l9��@�#��n�͂SV�U7er%�6���� �v�H��k_��v ȯ�/�����Y��7�K=����`J�v��y�wM���7K���I03G���H'������+T_a�x��e�07�jn���,~�N���x���o��n0G�M���k9�Z�o�p������R�����b�Fz���o����=�Hx/WQLN�>�@3v��#}W�Y:D�j����5�\�����?���w����M�I�O+G.?M�DlaA�6mJ��g�1��N�-�k3o�A1!�<m
�3���Ă}��\���g�М�c-YC;�=`��]�?�HJ�G�O1p3���/�(`����7�D~�ڠ�{t`#����	}[x�Q���p�Q�N�?�aN���t�v/|J&��+��� P�����U���:{�+��u:И�P!d�;Fi}
H���V�l�P�LG8�m�wg�|И�NR{�ߨ% 	:�9�~����n�����?P�r��J;6�w�*%�)C5�y�(�j��Z�+c�qA��vN����78п]G䓦7^���m;��b<x�G��k@�&�I��슡�Oa���`�ad"*���>���ۦ��=�d�s���?�RXD8���ܔ,"a���+"�56H��e�ġI���q��"�� >=T�(�_Z���	��{e[��L;f��� $��=�6ʚ��a5U�̷��u�Z����"�%O厥���C���� �;��9�6B�O���Ye�!��^�� lڞú4L�z{D��m5s��fE1�88�S�xY�j����^��E�%�8�y���Bnn�"df�%��Ų�NK�Ѻ���Fr�XP�GN��gktԅ,����JJ�D�� �`{X���E�7j�`��o� 9�u��J�C2h�j����4�eL�A�̊g��n �@�ђ��61�@^�^;1V&�f�5A���m�;�N�����p��~"�ۢfgK��J���M�R��S`�B4A)�G�sa0R�Խ+���-ʖU�.�*���|��|+�j��vwa-΄fo~��^����Δ�Zh_��wh��b���_�R��)��'H�{>����mvSg��>��-IɄ!�>,4��YY�KY�s��x8��I�����מƩ5�)������|��D���F��c�kjg<�x�����/A��
��&�~��(e��E��
��Y�|H�R*�������PWF�D��6��������v�:�rB��N~��+��ܔ��b�K�d6�H�X�A�Qiߣ+Kѐd��d������W�ſr�!����>��I���|�F�/A���i:c��d��.l�˓���ح���{5��8Rt_xV|V7��t�b�񷎰����t�k@ C�([C:/�K>�����G$J�;�E��%T��I���gd�*ѕ��
��n��YJ#�(�;�C��gS2(Ȣ�G91acF�sH�ս���[��q�^,>�=���0 ����M6'6�~|�Q웒c���wh&��QՈr��,�tv�E�{�#��r����R�$�I���H�9y���!��۾Z�.����VlO����a�rDɡ��
Ɩs�HSr��
c�r����Ȥ�=LO���.%���-�!ϻ�M?H*Z��7tƬ.�SжMM�%���*ͽnD�+��yt�1g���[�![������@��4��|�ݕPT��@�OdW����E�j�Ĭe�!.ї�7�(��GC/`��?C�L�)6���sLD���^���tXe��E��D��k7,_#��5����oAa	V\�L�75�}~}]F����*X�^u��3D�X���������_I���������Pmz�����i~�;rm�Q:�Q���Jdr�ef�}�ӶOM�`���Se
�-����ND�(�p����[�ٵ�8h/_�B�a����'&m�6�ㇹH�Z ) /3Z��̼1��]B�ğ�}�F�.M�Or�����^"�4�e��I���o#����Ӊ��FU���'xs;��˟-��-���o�'�K^���0�"����vL��@e&
���%��0B�r��6�2A�<�|�$K���]ێ�a�e)-֚E�e���ׄR?ߒ �����<K�%�~�m0kx�0�L��ճ=�]Y����;�t�OO�vx�HM������uH��+�,��=������恜�X�̄���>����ubu����~���r�`V�b*I}�8��ˏR{���=�������OS���+�9��Υg�;�I_7��
�-�w�N�?;�Z��W�y����о7/�u��j����p[���N�ȇ_��ȞKi���q�j�@�BhH�QX�ëm~����o�����1m�M	T�4$�+��L��I�r�>Yx'op��ݏGޑm����������ԛE���z�+52��,�\(b�SD��{�^֨��V���+��k�CJ~���� ���4��bн������4J�h�����o/ŗ^���3)�5(0m��.�	�pU�%��X�U�u&�� �R�^md #��9��d��O����*7G~?Ҫ��M�$!XT#;��9(�Y�D�m�6&�\�X�f���-˶�`�_@X�����v<2��� \
��x&��	��S>HT��������Zi�sˡ��o�5yb�ڻ_���N�������R�Spd�Ϫ�lD��-)�ϸ�k��?����Ʌ���X�Iw �C���G�Tԕ/d�}�>��0}������L���R��<�i�*�K���a�*+��jDú#�Q�t^�"fQL�?_��V|�~�K�-�*~.����W��,)�W��V �tN���H�{�����x-g�6�͈�=�r�*�ي0��R�e[�T�H`�Q>���f�r{����;�RbŌfc�G�Yq��Zˮ�Hx%���R�Fe�y�[���X�n����3�ꨔ6��7N���%�-���J�� Ϝ�_��)����qߪ��Dkܘ����;a}r��b�(�t��j�~��u��:t�
N�b�{�����v�B%C��:Ug����"ͷd�����A�X\�W5��, �|	����ȡD+��(5�̡�_U`u%g�+>j�8�&��T��k�^s����A�{�fi�4 v�$�����l����w�QxɃ��N���Sr��g+�e�.�^��5��92��D%ꇤVg�U����)po�_��u)m�D�ê�3�'0[_�k�A��B���c�T
���?v��������ȤW��ګ�UW�L�Ҙ~���x�e4!�m�
�oFP���0�l��cJ^ܝ��.Y�Ɉ{e�[l�%������N��;����M{��ҞcZ��g����Zu#����|��T{��5B8�}��FJl�a��*��A>�0}Ҕhd�p;x�F�`�1��KrBc=��n�L/�kP+t6fAږ q�l>�ƛ�v�޹.讆�=�2�Z�2���3�W]0����փ�O�p��GY��g)#`A�w��F*��k~���ݯ�7��ZM����q�� '���5�M��r��KR�<԰�#4nRK�:�r���p�j�����F��������_I�KD�;�U�c�b^�qOY��;۾��9'v�?�����a����Kϣ��7���r3��!����\=���)��Q)�P��X�Mu��L�ֿ���DL�_��:Ul��#4�
%�:=���Ӡ-�P���������#\��3mj�W�m91�Q����� R�ɭ�0��N�|�84����d���ae�Ä�q=@�c�]�xNArh��v'�\Śl��3��!� ���%q�@�]��׷��gO�#ah�SD�M��8�k'�9���2�i��L�nŮj|��*Jb�kj=c����G��@��k }�����ק��~�Q���"����ݷ�ה��!8�񳅆��ND*m&�eTz�q�N���2a��p[�F6�;b����_ݸ�]Z��yOʔQA�Ʊq���zd�~LFX[	�0�J��M�W��5`��b�a�G5Dt`V���]�Kd�Rn�/��K6���� N��^�?Ov 0Y�������Е(��0H`1�%D:�~�Ų� �Ÿ^��(��`����H�ȍ���E6^|�fu�,�b��u�66��0��(0�~=���eP�*�5([�S���h�]�hU����*�X#ϾЛ�)�dN#�:�����09���D�-���Mz�+�(ɳ����K6��)7����;	��t��v�8VɦƫL�Q��p܂�N�%d�_���-�ڙ�e���+�e�Pd2�V��-!ޞ�p���~c��Y&�'in���q������gO���V�$�F�/=d3݂���؇4�G�#aM�Uن�}ǪYYB޼/ܮi����Y�tjORƹ�S�>;4���$~��3���?63����|�37B���:�}*T�k1�0ʤ?��@�|�v[�?��^G�Qh�@U��4�(V�4̴�{�[�|C�[JkWx�e��|mD�AR)g��
��Nd����.�D�++��h��q�8��0���$���VљՂ\L��g��k�����#�ڢ�W��-x�n%s���^�_x�zb�1�Nn�IW?���/��av,�C/@�<mA'j�T�C�^ZkXF��t�0��w�O}Jx�0��r[%���4����
g"w�ҵ��t�^U�aJ�>=ۺ�u��,����+)Kª�(�Z'{?x�oUZ��i�OOĪ��ȼ$",ϱ�'�Sء�#D�}lWӪ�	��`_������M����Q�Ԭ,I��kĠ��<n4r��\�B������*��w���1�e�-x>��2!�9���wpۚ�|���/p��@��� ��,���#��z̈9�
'ɩbn(��yJ�5T
҃��Rw���&(�dL'�d�ʚ�����Yχ�V��wLNu+�Մ���0�1���6#�	{��NS�3g�fT����0UO
p����.܅6�L� ���o�z};9� |!���Wϫ�`��t����e`?�߃�}G��#�2	�������X0���)�Hq���#���q�!��.j���?��9W��$���J5� R�'4�z���ޜX 5$y&�L�U��mv�=j�\"cv�z�T�1�"�w���鳑�H���܇�'Q!Z
�>��ױ����j���K�4�ϋv>��-iw�g>�ʾP�e\�2�*������}l�K��U�.sh#����A�8����X��aі�Ѫ��SU/�S���Wh�A6:$j`���IQ�o4���������+9`�ԍ,H�M�;*=/#8z���2ߍ��FXR�
�J�8��J��ID}�����/�׻xl�Aj���\[ܒ�A��2�eｄ���A4CF�.<c�XMp�덍h�6��G7�\p��&��F{�|P���gJꠈ�H5�l�_�o���}Z�*1�x���O��u�����������ұ�ä�*�o��ǸP� �k?�iu��3Oq�کn��n�_���UBLe�)��K��Q#�(��<�+P��1���6�����*��Ј+���G�:�秞�@��6��@f��ܠU?���x�l�EA�_%2	U�����������`˯�|A'${OT�s\SaV��U��絞9�����<��$�^���v|6
W�l �%Rw]>.�1�K���4�H�\pCq���B�.B��Xp0�o\t�����Gu�p��%��C[Ǝy���,ZҳC_�"����pʦ6/�V��k���
�SM�I�ndE�T�U�ڄP�h�W��N�W^��}���U Ø�W���-١$:�	��U������n�!8��r@�����:|�h�?��-��VX@¿]>6����6B􋺾���SG�q��M�x^5���Ǜ��Z����/*�r�yru-��������[>�]�B�(��������H��ڛi���F���]7}G�;|����!�|U/@�,�GG�ӎs]����:�nQ��Eu�)�]`i5A.�Z��ۺ�p�n �q��y �k"�/��}UĨ"]\�ͼGK뽋s�%�X>��':B��e��;��Q�H���Pc���BPJ��`�<�Iz撿Q%E��`���N|���&��:��ӯ.@z�F�����+ﵰ�lx[=)�vSZ���	�uE�2k���zkK�+б��5_��xj�<μ��>�W-"��*S+0E�@O�\Y�	�G^<�p�娳}�S(����� ;�������˗�t��?�u8@m��(v5�VVV�$�a�ms,|_�ŕ�Y�|�#��>G<օ*ٕ���`ϊqN��R�+0�d+8B��KZ@Mf�Uk!��~���蛻l�W�7��oU{��ļ�8g+1�:T{����"�%��,8�7�Z�|Bp��A8�/Z�G��CP��ZaD7���-� j���-lm��e�Z�+t<�8e��W�h��{ �F2�\��`�͊׫1$]=���'�+��>b�����P� �󫋭$w5�xe2�2Q0���դ\�}.�$ڡc���]Apo����$����eF��T�E#iʟ�{�2a�y @�"�?�� Ο����V���͘%d��,|�l��$��p��(��U^��-�Y�/����q���e�v�zn�2O}+x��s�FWWu�Ȟ��7��P�^-)S=�0(ĳ[;$��z$�=�%1�qCq"�T��;V?k�/|���jܡ
w�P�*x�֦̂sEƕ�ank�Q�^[i��gkM�0��s�ɣ~��PnBGMb�G.��qiK�Y�����D�K�^?�t?��?�|m��M��֠ ���|C2K��?�����;��1@M��p.��[��`J�D�Į���;�z��Yc��֪@����R�N�|�5Ŕ|C��R����B��o�f=2�^2`|_O��Ҋ�%l��O����*�ް�ڿ��q�����;�F|Sr���h�^�0:���ܥ{���x������}�	KY�T��܅�&q�q�ѓ�=�(��
���z� �[�0.�����,��U��~��-!���C����!��B�~�Ť��nq�YHW
P��#b|�Ȥ9��2���CP��#�r �����/֕�J����*�����\UUBS�`e>��LoRF�^�����p�ۆ�J��"�3*�Nr��n%w�������w�g�+��i�������z_����V�r�Y���/��Sn�4��b�%;�)��x��R��*xMxkw� T���'�\?6�����+P<��h�f�������_̋D>E�����j����0�q��K�������@�Bv��~!�^8�`�z
���]�?&{\Ͼ�[~��`�x^|ೂD����R�D�̑����ǋ��lmSf,�CJ���b��YX���Բ�#�i�뛋@�$���ؙ���z;�%?$� K�{��5����?�W�A��4��ge�L�5�O�fb���4�8�;a��Ar��΁��YU�ԕ����?B<�>tZ䛺����4a�Pcv4ƕ�|)Y�P��Z�`�"��G��Zbj�9��Mұ��D�<W�D���P�������KX~�i��D���?�H`*�4�����;���	3�.i��d��c͂���5 
i;�5�1U���([���QϨ�s[+'�}�9&��2C�z9G�z��g�ʸ쯕�G'W\��Ù���֐h���f�p�Z����E��j��o�9�����Uj_���%x� 󦷤��_,�@lG�-�CP���bzᜨ1C���vk���y\?�l���+蕪nMOӎ>����rLȟ
�HI=�4@�%����&��8�	�"� .�R���T�c�'Aѯaf�:!�.����f4�dQ�Z�ϊV��z���6�
:�"���L�t�)�,�dh���E[�Ze}ݒ��S�]��mП�w��F����L��.xm��ʞ7�����z<@�^$kbs��oO�`<�;�7��z���|*�* �V+�H�Ѩ�|l%Zp��
9�y�l�Q�RÝ�A�b�b�m5ǂ���f2LMD����hn��l���Ӭ��z�}k�l��GT[��8z��>��`n��w�\���a&� �ߨ���u��Bވ`�l��=
_;iM˘
�l�Ƴ��ʙ�曅ۊ�����1	��MDv��0)�����yɉ���
�
ߪ�Vla�?���1�bJ�8}��ƊD���
��N*��->풮����oǘ:�A�L��ȭ1iv��� !Osc����9�63=��Y��P��T2�����ƔM�֊���:�����^��V��ׯ�<u�K�SL�H��<�����\��{���C��J�˸�z�專k���rr�qAu̕�弅��օ��!'r���?j8�A":��Xk̇�/��j\�ji����>�\,'�n&X� q+�z��\T��Ș��O�uJby����]�;"u�P� ���Qm�X�	��{5,d~�F�z8���j=O|S\��"�}�Qb���ޭ3<����ə��F���@;�����Rd��^U���E�t%ɛ�=?�RP�1�Vs)y��n>|&��U��)���� q~*�yv�@���v�*a����ĮJ������� �m�qX,�S\tP&f�Q��8�"1��w����R`��ݳ��`3&ļ�\�q���i��62�����!���ױ�����+x� ^c���B6`Ե�dĤ�����P[��8 !��ߺW�x"���ib�ҹA��gjB�nr��,�H���3;�R,�������^��y�о�[��)�>�u�c�sI�3ꙫ�����*�k��z�K_5t}�b�e��9/��#ک߯�A�6�}PExl�Ǎ� D�(7��v6O�.�o�SZ^��g��k�ۿ8��l�)�G	uT�V�i[s�,i�x���~��ؓ�p���� ���qV4B>S�ۥ�;B�w*���<8����M�(�Ai��Jm'6=��[�>j,$������Z�Q���23���f��J��|t*��-Px/��s(1D.��Si�e���X���sc+��r��*h4���[��'��|���*f��9S��	]l:��}�'
5��~{z�O��_Ŀ}	s~�;��f��=q�2���B�(���c���ҹ&Y��z�N���of8V�ߜ�Z"z��'�̋Pd�`%r����)c�Y9E�2������&8a/0��G��Ӣ9��B|Nrx͸5N=��т\��my`U_K/Y���-�ː�!7B����5Y��0Σ��]�E@d��a��_WI�����3�3�z^y���BX��� ���
��8#�Sg��n4*N!ۦ�AIsf;i�'���j��PJ}������O�o鱠o��␼Q��J��f��V}J�]�i#Tn?�Ӓ��W����h:n��E����yǶ��z�$]?��;he"5V��+C���@��#kz��ۮv�8�t ����3g�.�ղ�	[��73�!����b��5�����L,()ӉL�}�iD����V~̵�ToT�9ظWm��K�F����8Sl��=��mڧF{�誼U�띯��Mm�-�OwC[��9���f/��� <�#�5uFο���K�y)�N{���bۯ7����,�@�1R}c�����M��Y�dɞްxh��{Ϫ���_!���Z���2�k`׺�������Ď�B谿�9�Ѵml���\�U�kRU�vp57�J���I'��C^���;���%[=>�;�Vs����Z|��>5
^7����0r�Z���HQ0I��=qkAC�v�t4�z�'���cs�v�"��(�r�:��76cd]������a�1)V�Kq�U��Uv��m�F �#ƴ
̏#k�/Z�`�A^�2���m�,�����n�.�_>Xv�E�����,B����b�X��A��!�{���+�u��Ɖ�
yl����E� з���Ot�!��ք�R�#���w�=�gVd�k���⡷S�g�5��Zجz�4������"��p�{�iM��w#�tz����*.��*��<;�2�/Q	⍖��c���G�3�m3C�j!�b�33�{�]d�O>�y�ZI����s34Ң��tS0ܟ{钄!騕���p�]D2���<�4s���ӥ�s)�+��O�l!�8�-�p���K��T�4*��7�R��#��N_��Y�Z��+}J��_�����&zp9���*�;��x���U�Íl �����ײtu���X+<�e.�p �ѡ�Zh��``������u~cC�Dh���Y�9�+<g��T�CC^u����&�������q2t7ӧ��K]��O�%��J��ڋn?�~�0P(gq%+(cV�6�G���&iL�/(�E��Wħ�����K�l��Cֱ6A�]C�u�=�"f	�"�����Ź����`�'F�'�U�CXZ����=����fn���L����Mg4�2 �]�M��A��H��U�vb¶o�qw}z�[������/Pm��/\�w��KD��h��
���$��9ΰ����&�Q�M�%>'I���j����cMX�⑈�U;\{ NG5X���
�bV�&,+���z�?2��g���C��?�gM���i��rH�L5����ꐒ`م����ރ[��͹�Ц.�	(��N��y)��o�,���������A95��<�Z�Ñ�)RT��$>����^�9�6�SLi&Fy-���r&����,F����kq��Bv��!EϦ�V��>�e���(O�->[m
ib>��J�?��L� ��!�bfC5~Y���%$�#o]�-�UP�^����,yҕ�G��%��	0ED�t]�f��xF	�1r�Z1�(�'�7f�4E�P�^l{${pA�><p�,�@qDr�F��"X('AZ)7�@&����Bmی�j(otu������A�f����T��+jBYl�׹F:�oom����Ӆ��~s81���x347�u��'y�����D$(x|^��_#�4o�ଦ�-��2���������Y�0�(H���lQ�*�Ą)�,�߰���cvV�
�VS�{n���9�*R���i�w���'-�Mƻ y�e����o�f-�մO�D
���PvY|�V�� -r���c�E�8LG^3�Y�%���l���/u�M'�C=���=���j����4C��M̃�l��V�ueXϢ�LSK��&k��ɍ�
��}�b ���w��fSg��TV'� 9��&�z����У6\�^�\���,��C��[c�	�5 ���T�	����n_�*>�܌�҆Jx��1�6~Bu����!R�|��6� �P��)��ld+^ns{�#��!;"+�-3����2��F!���6�t�ӎdz���ǖ���&���5מ�[٭�<sĂIsN�v�`�'WU��pj�P���9yJm>*?I��n��:�� �7ͼ
��3;�e�0�2�2(��1��߻��p�i�8.���K�L}�F�����I�쫃f���vd�Lmuwi���,H��RN/@�#G�W����̍����"WZ����_�N29imlKC�c���9i֏[����|�z`ů]����Ӛ"i����3�q8,h�=��6	;���>j�Kr���d���ͩ�TM�d	s�2�*�*��[N{X�'�c�M��T��4����}���)u�� g�M��<�dy-���M��kHo� XT:Vk��B������$�]'�[S}�c�MPo))�d�dZ���̓�}�Ԙ��lt&'�6oȆyn�C�&�o`�@,�;G=6���:׮��:G�)ҳ��sx� ��v	
�^�ِ����t�i�7GV�9�D@�-v�����c���4��l�(1w�
��NPϫ�-������ �7�S?"�-@��鄦sѨ��=�b�]Vr7�EֆV|,��-yg�{�O�)s9S�d}�i��ED�X�^&M�-52����K�������M��{#�	�e�fR�P��t��0f�t���o�<a%D��,�*�}q�"��Cu!����Ｉ:��-y?oTp�k�B�h#��0��rǷ��|�<dp`(W�Y#М$����&���Y[N����4pW��a�K�ڪ�J�.痶h��s������G]��盰��\�nO�l��=P ���;$��ԍˊ7u���⼢������/��������o ��`ɡoUH�H�� ��	s���hĀƆ��%k�Jz��Bue=��k1xs%m������n��n'�;vոi�a�s��'�ݎ���}��4�"� �n��=,�*�fd?	S<��f-�A�a$'N�nYZ:a�����+׿��̼`�H[}[=���)3�7�7T������f���a�#Z������8�>o`���!6B&�WY������ zZ���N��N5�kǛWҊ���]ʗ�޴�Au�B�n��+�jש~qhU�������v��jqk�x�'C���UY��~$ �Z'��$�ĔR�%�]
�t&.�IA��`�~��H5�>�Nl���HMu��j��nO��8��4�2[�9��~�T�Ľ�����ZZ/�@�a���6Ҵ����t�0&�O�"x���O�NoZ��f,�����9�j�uT:���P��F&�b�"����:�+
S�z/����<���Ȟ���>Q���bh��R�VTs?p϶�z��ݱO�'���^���$4}�i6�m�}[���ԕ2�}��T��d=<��SVB0˘L��q1#�z�"[��n��[�)�@�S���yc��o������bC:ޝ��N|	<�����O���ݟ!M�`_���2�p�ue�`�����~A�$`�4��j�9!%�������TP�i�:�d��+(�����Q��7�LΦ��ao��*��}C|[8����ǂ��)�	b�8ԛ���z��:0�1��������ܥ(,�`X2�$�[��0[��2���D^��&K,�bt�d�� ���VS�*�62���U:�zr�aSG�{��5g�x�Ia��r��њ�%�Kv�/QXao{��3s���.a��l��o��j�z�<1�M/X�Y�U2V��zFRo��ɴ	��t����
��o*�D�E��e1��~��M�<f*���]V�yHdTN~=���<�p�	�`�0</u�b�+������Q>�U�ch�4G�Q�S�]_�NYF>�M��`�Z�f.A3z2<D���5�dխia�Jn�}�P3��5mbc��9Fߓ�8{�2�m��}"X5@���=o��:���yt�M{qhZ��`{u�Zd��>�9%y�;\�e�*��p�I�Y�m|֜^��N'�t�d��ݢ-E,��R�0"��X'6�ϡX�Fm{�E�K��fF*�3a���~�Wr*�L���]�qpR�"N���[(�\[2ٙ1����\,i�@�sE��֕�̠Ҹ&��e�C��H��Q]t�b;ۃ?6n9�E��3���Ҥ	�?���Sը�S.�C��hb@���<���K�Z�%{����Yjm�S]B���֐�Hw}�Ǳ��ih�mk��Q��\���P������Չ�4Դ-��}!b��q���Y_+�`D��<PEAI�:�@�ҏ�o<�S�_Ŵ��K���CQP4��̐�X�>�Գ��(p9�T��3!Q���ߑ����H�M9���0�I��|y�3�C���a�k�ȫ��GP�|#bS�y%Ů�~'�/�!ȭC�1���0d�Z5���d�

 5�5Qt��}F�\�[y��YNlQ�I�u�6omd٪�9A�=�����5]�'���c�� ��cY@c�n�q��٫��cX��\�Z�L b�JD�����X��#9$l3�Ww�'�V�=�U�m���=m�H�A؆r:վ�U�=(��t��/��Ŋ�_+��!����rif����� K@B`#����u-�����Hwt��b�g�
�{Q�x4��9YB�\��r��-�6}��Wf�w{��w���V�(#��������<����[x���&��r�l���
�ߥ��Rl3Rn#����KqO���Fhc�����lgkE�RM���Ҹc�?*;,���+��JV��X�I�'��;��ؠ(a�܁
9~]NT�hܷ�2��1�����4ߙ�A0��� �ϖ��ٟ�k�VVb��7�0#�� <#%c��	\�B��@4)�cFY����-�������+���qAw	|v��$�w��g��D%��y��)��X��3g,��u�vv#��(���6w'��Wil�o�7�Cg��;<7(4��b:� �V��8�������7�羇�{k��;��ϏE�!��0�vX\�(�����`c.Ν�Y�v�X��4����]a[��t��1��TL�������pR[�PT���[&ˬ��_BA�f($C�=��m��#��q��E�;Z��(��{�IeWE�B�l�`,��1��<X/�mɜhk }�+% ˞u� �DNUe�%��iE�-u)�ֱ'�Ǿ�Ĝ�Ӕ��;��.�o��R�,6
f��dޡ���XK�dHM\1��J���A��6��3҉t���jr�2߾���,Y^��jv�X�i�P����H�e�G!�`L�V(XZNGKO񉮬���K�Ҩ�Ӆ��)F��ǲ��fn
�>�5�E��*���40��Oy�LEj��+��
͗��4v]j��JԪ���tE[�M�z���U�<e qM�*u,�&^ŪO��L=�&NX#��m/G9n)%��n�w���K��<�&.A�'&p'��/���z��nQ������<�~+4I(��,�e/qHf9��k��Ѭ���@<�3��Q�#臡�����{�c퓯�zl�<�6���*�S�^���g�%Hy`(g�kd]�u�F�@�������.,>%���"l�	G�︋�G���gh{'�/��s$7���I*��ҟR"�Ш�ھv�j �<QH��e�/�W�t��d�����㐹��'Z���G�_o(� ɀ>����)�8�'�*ޮ�dUy���}>��ֵz����s-�J@�Cf�+@�5Lճ7��F���C��d��5t�&ŷ��žѓOH�b�	j�&�P�c�65��F��,��Rzx�ƭ���
 +ٗڼ��G���� ��6��g5&M�a%h���#A�����inT�h�7O��kl&����s���v�Sz���"_��_�~�ZP�� �"�5Bur��P��c�z%����;���P\ء��Z�(J���g��ۆ����h��*g�D�����A�M��=�h9���d���c����nr�w3�d�>��!�/C>5֍��KT;n��FZ+����{�<V������7-W�J/��[`��F���J�T���]�ﻓƏ=X��{L���O�Æ��C����0Kl<=ƾ�Ym��?(�w$�CM�h����������[� ��X��Ս�0�L�La����ո��ZQ��%�dDmmv��V<��zo����q��&��W�����W��S��^�hc28�s�+p�=��P�>yW[���1�����sބ�{)p�Y��C޳2Or����wrVca��Qu�)�l�R2f��T{ ������vk�uT&�s&Obg% l��Y��4����4nfp�#5�Q5���n�d֤�ެwrg���F���$�C��ʳ����Cot��+٦@��8	���,ӿ!��Yח�����v�x�uR݀7]�ߋ�I���8�,)��
�� ��\���녈$�]1�/��-L&A".!-"��V�YS�Xw��/d��&�kpʛ�h[�V�R3C���o�B�sn�ũ��@'�����o�A�:V�y(�HjEtZ�,�y�Ui����N?��) �^��e���Vw���Z����7����M�#-�Z�#O�����p����oox��d��86�$>�G?l��b�@I�,�7���AOe�٫ø.&£٘��h{�1ٗ����(��T�������e.�hUQ�O|�0��7�W�:��n��y���O~^�\��vO�g��)���U*nH�8��2az�u;���%���O��{P����FB���e贺E�(���bOu���^>��x�ٵ�{(G�}(�V�\
ﭣ�fI��B�d��m]0�^!@*�����rE�[_����@o�_Vi}y����<�;=�rF^��a��ԁZk�;u�r�P���Ñ]	�q�ׂ_)�t���>�2�+/i��Y_�=�B�Tu}��WuHT2Q�`}h�YRG(|�tLl��z}0fr�׃��߉^6<�KG:ǗӔ�5A
-pfX��9�_D�?��Gs2��G��'YC^{>�P�����%*�YT:�F��[n�?�����x8�����]���^31c�( ��>�ܖ-��OG�~�fK��y��Dr�ۍNT6!u��"��/֚��U�̀���r�^�LL�rq�3�0�8_;�5�3��l*ZѮc!f~x��]��ehzU�!Ƅ���F|d��f�J�j�Y�3h�qB5����% ����}џ��s�V)�D�9�^ 2FS�Z�:�������6R(����a$|Kw`#��|!$oJ�J�,�"��3t�8xx���z�%�ᨾ���L��G�+KnC�ް̉sG��
��� 9��]� �
��B3�pz ��`�p�gi�������}'���54���V�'�jW�0�j���
]ӡ��L���=t.W6�ԢWM>�%�k�F�k}�J�� ;c��3VA��ֹ����ظN6R���0����>L}SM������Q�n�W9�S�|�<[3X���U�?�T]�:Ts���7��H��].��1�Y�	r���^i�
;kEbA��A:{�Z��<��S��}�� z��t�����&r�
շjy�U��"b�;%�=�D�XX|�V��% .�*�Z��H�$_��	:�/�2~�����'��q�"��u���"��?�!�PVW�s~�p��g�:��˴������VG���!0����4��/l��d�g+�r�m{��t��w��N�hQah��h��͝�!��gfˏ�Pj-��������#˝�˕S��C�&*���d�I���(۟sBu���
Ց調4S�=Y�m<�_Pho�I��~8��7 �~,k���t��=��)P:.k9���-�R�'�-�a��SL*(i/S�M����B
����
�Fu%�W����*Cd�Q ��Frή�B�!�r!Z� ѕ�]�:��;F�S<F�,J2uM�⢫�7�;���|����eVO���|��q>9%�@0fi��|p�U��*��Z�'yI��-BD�(�8ۤ�J'���L�������҂��A�����$��m���?��уkI�.�c��\>�i<j�����`��+��y�e�f�V��eR��2�>d��3Aw�'~!�	��|��C(��3V�E�CA�U�\�RS���ջO��&o䁾t���R;�R6]H*����@�:MC��*�gu�E���u;�Q:��dK}I&Dbq��:��N���ϵ�h�Z6&�O�{@ûX�����Al8�=	���g���!7&�,:�wq4!̈ɂ_�U�BF��W�m���C!�Fw^!5_l���g�u�h~Y���!x�LY{1�!�{eų_�l/�L�t���W'=���
��߯V��E��Y�.a Dޠgmܖ�6ˀ�}Cw�������.��'w�E��;�L�-O�-��?�J%舯Sݰ�yYH^1�j��mk�E �9p��e�<���>ݥ/��͂��c���d�h^ݠ7��{~���_�@��O7�j�iT��
7��L�n�}�*�K+4e��1h�N�͡��=}�Tߢ���|K�^�էQ p�B>�}l�p�zE�J����q��-�Z���p0�A(�߻�Ł��H�U@]"�ݺ��FW"v;�mT'%d&��s3�<D�k�M�VD�G���r.P�8G]�*�9lT�������֛��'m�-h'yp����"7ޚ���A���%Vnb{X��H'&��yc�L+9�?� �Ğ�X�hr��>�#� ej�y��憆�=*@ݥtC�
�}������9�YЯ���B��EQ���L;����gc���*�K|(��m�=���Z��e�lr����SA��p��pٶ�/S�0��sV�Eα��D��_u�ͤO�	�wF�9�:�\\ܩ˓�͵����������+���1�c�lf'�OQȭO�`.�L1��>~��	������L�z)CO��p;�*�ʦ<��̼5�� ��5��)2��&R�l�E�
��7_!IC��>�4���}Q����-!!]�wp�w"<Ϋ�	P ��
�P�h;��$�IW	|h%�iB�t��X�+�/g�=����yb<V�
ay����x9\=��&��<DX�ZT,��'�����´��X]s&`��"B$�	�i<�W��D-��ǤR��/��&A�� �J�D&��;p/���Ai.���t�YK`ps�7V*���,�/C�w�����ڣTs�ӑ6�+�����@�-�׀�_#�J��A�gԳ����{�&��I�` �J��)vVt	 CȌ��y��}�C5�v�:���&e��L}�-�m�o�3�g�ڎ=K5<B�\����+��e�N{\e���o����YN�	�h�'��l����_m�]�{�`e���h��>�s;��������%0�%#�}0i�K��E���B�(݅7A�xc�,�I��F�U*�L��ㅆ&��)����ܖ:�0]����8�v�韴}߀�;�����y�����r�[�"�袯�V�"���)י�B���V[`�`�@������=3y2K˹�UK0��uC=��^���sF�����H�!��$8���� a���B"��)h�#d<�����A�BGƼ�e��{�!lt�ِ�XM�ذ]�ZI+w�']Ψ�#�OCb�pZϚIy���G��e#Q�.��0-TcW��B��s����%�2u2�CfpL7C,���(�"K=xs'G!��??:�ƺ�H�^�����R�@�-�X�D4��B���C<���C��p�CJ4�G���}�?mH22a�����cD��xn���R��)�����(>��CL[y�_��u/����h�R�*T�$CA��-�R�j�f�R�Ե�����% g��.&X�zB:����˱G3cn�p�u����7�U��H��(D��+��B��y ��ۺ@0fi,� X�����P1�����O��1]�֝��ε�u'���6��K�W_��o\D�M|�6Q��ql�D7��H
��F��B�/a�wG����B�� ��O9����ao%�Q�Pq�9t蕅(���F��jΝ���Դ��Z�x�go2�I��2�rY�!�Ov���� |{���[`�K%5�Bx��3#���\�>}_h�<�r�
Ss�E�v.yph��S����z\!��̑D`5^�/�1	*�����ȩG��7���{G�]|1=�	~G��&��_d����A��Z�N�L�V�w�?�\��g7n�SJ�oK�c6�y�G-m�uj��U�2V���m�������R�㣦�W��3�is>�yI������Oӄ�����Z�n����9�jc���[k�]�Xn�7����hT���Gt��r�>�ԟtNz��s�|R$H�hإ>e/��fvo��=������A�(q�Vp��%��a����4�{/���k��B��CG�	nW�&�d4�bՄl��5lLL/k����j�`�������z{�\����b'��cJrG��7��Կ���`�y|hp�"��]D�Ҳ�>��r���o7���.:��2ހ_�EUK��hhU=]�6��
�Bc~��j�1(r�F�_�'�K�?�Op��������g�ɧHL���,|Cb������C�?wkXڔ�A��:͌������F���>�F����z�ٱ��knrZ��ǒD�(S�HD�n��է'?Mßl,#�9�+�q��f+��~��_,�ϩ���?1ԁ� ږ2��7�jsڏA�q�-�Ge=Z��3��;`���Ot����m��*WHe�&��e��d��v��x�.����Az�nj�)��@�ϓ|p��'�+b�d�½��X&d��0|������]
�u##��-��b�u܏��Zy��8�n�W�K�?�>��t�X�~�*�u����s	":ԵO�(�v6��<~$�m�}��[��*������BB>�Ă9#���h��m�E���!��UO%&�Zɒ[��M&���L�m��1u#v��S���$.��"�p�5F�Br���ob��Ym�-�a����Y�d�?���	��4wB=Zʓ��:ܛ����Y]��_f��9菶Ӹct��gS����}�h}8�E.5��I'�����
?� Hބ�%�fj�=M#�)�&����T�M�a؆�D�	W����H���cQ�"��uD�*��^^k�$C�b�z=BD�������N�	�;�HE`>���=paz��H��Čd-R��BW�LH�@��%6��b��-g�� G8>h�¼pؼT��b{�J�\���O�O�v嶻E�>_���x �[c�*Ǆ��!�y�����^D�T祱�.��ad��H�<w��ƮԁS~��#���wXs�S��?��jx�.����qf���F�g]c�).����;̈́b�-�E�B���^Sq��­���<o�`���~�D���h����ޘ~sk�N7�e�f�pH�ݞ3�Z��R[c��v�z�帩s������]L��h�����GQ4��N�@�?��*U��~���!{F�U�s81�{�wF"E(�r��m��L�'g;/�y�Q�,1
n���6.hy�b��(�.��Yk����r>p�a�ڑ5C������fU+�{�!�	�cn�HI�})i
�t���x�%��E͠���[_��{�7��k.��bg�H*�����2���`�n�,Ȃ"�vO��l<�hC�8@Ļ�]n
�V�%����󤠸�RѪuGb��7�uMd��w���03ZS�B�W�0�9���ڋ��_Px����yg�=K(U��Bn�4�H�Qu9�eڒ⌼��>��4�mEh�����B&��v2\όaq�E�.�gF՟��%}���F6y�~f�F�L�N��"%�w
)J�n��*V����Ff�*ވ`%o�O@W0Y���| ~ޙ
���S��s|J[l����)��S���He]�ѹh-�&�n�r�jupIRN��A������KO����)�L��lď��̿ ����&�p(�a_^Xd������N��<سw {�Ge�.q,��IpX��>�B�eZ��� ��JJi��$3�5M��/�@gs�bu/��>�f�l!)+��QbK\��y�ezŠ�5�giq��K�(��~�f����]���a�]��N�ۧj̲I�t�e *]�HާUV���jP�
O�f����Ԯ���x⹙�c���V����hԮ������P��`�VA6������f5F�'Mzmπ�dr�%h=��� �9kO�����@3My%�z�^�R:�5TAx�;���F�`_xˏq��Y/�U�$��N��f��(�T���;��q�|���5��0�OC�>�_��8bx����
����t���#B}4�,�ѝY����ܛ�'Ĺ ��o��$���O2�,O.V�J�L����+�H��^�/=��P(��'6��H��|�/�rQc5wLu�#����%�M:!��16~XN����Ǚ���Jq�9�c�=�a�@
�'Lu?�l���m���o%�R�u���H���_�l5D�Do��h3�s^|�ͷ{Q�*Ew�B����܂�a�[G���ަ��y�z�r~]��Y2��m��b���&�@�]��C-�W��]�!:u|Uxy?o�l|p�`ShG�<o�ভ��sD�;���a�Q^f�{dP�#�s
�4���g�k[��eP�\wE�A(@Z���4���_�ꛂ>��v�X7H�_Ơ�t�wH�s��:;����t���3J�����C��z��9�b�	�m1���VtPs�.�w�{�HKz��55H�>y�[-妹���W�7�ss*�4����)�y�(|�s�8uS�i �����y=1-1'k$]�>��:ke�����?
�%���C�?^�o����8�3�n��sM!��0�i��oQ���콮pM����twT��VhW��5j��L�1��Iw13p�eL5YW��t��� ��j����a+�X�%���{`�bG^l����J�Ǆ�h#���3B�Ξ��@�s����ةp)�{o��1m7L��'��2*$���*����_���(o�]�����o6�x+�?��6'"�r���H����˘塶I(��h�=\	RoOX�t��Ǫ�D��H������a8˓���6�#>d��*�}ɇ|+r.tW��%��iY�dW$��Ww�k׺I�����S;-�Eh�`3������zKɣ7i>�h2�@����A��ޅ��D�m�<���Ƹ:�D��;L���tT� ~�A�X0��3�h�M�R8\� St���;�m�/���ٽk?�.#aK�m��0�.�f4%񻒤���	w��Y�#�4�|�-x1���b���)�%h��ܮ������^��eH�u#n)�R��-���S�d?���e+�%��e�0������ө+'��f�p����Sj�w����Kyv�?�H�f�[���p뙺|n�ϊ��E��,���ĮH[�AɄ��E%��y��X�n�h&qT���" �.;,�#��yK�<w�զ�xJC���]�ֱe:�������v{���:<_���"�Gp���χ�xF��ܓ��A`��JPN[MXi�ۂ�ٺY�9�x#ů�~��UO��H�^���t��^ڧ�d��<ٸ%���zu�Ļ�a����z�~r����-LhX��L���k��e�������\ԛ�}�u�����Ҳ_�M0;+4��e��`�l� Y��XHiw0�����B����������N�K�lM$��{=�s���h�M��T�&vk���"��ێ�JJ��G������r��+�# �
f9,��=��t�ϪwV�^�dB���o	���Ygu?��=��x�q���f�*��D���<^��Dlm��NKJ�����m�Ҡo}��B};F�mT�G<T��Γ���l�,�|�By�D��Y�U��s����cE���?��m��%^U2˧����I9�N?��5Y9��?�y��ڭ��<�ƅ���ƅ�����eA�����w�4��: NnR��J�.�X���g:z��j�.�*a�_S��2�j��� �=�lS��/�\�s�/�|������:��YN��q��,�o^�	��9$�u^l��tt����!��q�'�Fn����S��D���l�����"�_��y��$��724=��KFc�if��o7;�DɁֈ������!!�)j|�i��z��$^�Ƿ�>׍�cƵ�B��4ϸO0�J�>��˻�q{Z�/���@U�����X2�qB3�h��V�wz��f�=���ηP �F��1z��[|H���-�tR�w���>y����������ۛ��e9��z�3���̊$uҊ� )3��4��3�$ 寛�q"!U$����{f}:�(�������
}����,�C�nP#�Y�� %Q�Q��+.Հ��P�GN']�W7���
-\����\ILm�/%Ħ�� �x/�6#{K�񿁾=���g�4��������ڱHZ�������#����]�9��1��'r�,����bȿ3=���� ��'C�g��i��;g�>w#F��ob�|���)�~[Odd5������\��3w�M '�|�����]���h'U��I ����>җ����tp�����)G(&����"	���R�ckϥ��/��p������_�0�}%�p�u�v��}7؋��N�;���t*\���`8(L<7���	�"O0�YK�*���t>��w�(4l��|�ewD��g�D���v�m���o6��wɮޑXŸ�	2:@���v�*��m�%�AA��4�ܘ�>�ۨ�Sb����?G�Ö�����H��+V9o��W`H�06�ց�	����Vȑm��`���������ݲ��G����5B9{���J�����T�#q�&���nn�qg�D<�b=�0��o���R����x*t�;̔�Nny�R��<r.D���`c�	.�߉I�|��!����@\^Ot�>K��,�8>�Xp0Sy�_�'bs�s�gH�,J݇�̯{�v�����CV�*b���;vĆs5�ҋ�a�,�ʒ�=趾��ͻni��'
=����ϓ�Ѹ�����\�?p|���F��elG 43��}�ǂ�R&�当K��NGɄM�zG�;ՉY&�u��K�����yvߐ��afu~�5o�.�qV~D	h�MT$#-g\�6w��L��:ԇB�nYO�I8Y��i��z dlNp@K{ ��'�e�ݻ%�:4�)k_�9��p�X��mU����Ө�Y�VN��/]f!���g�2eQ �BJ.�h6'������Эl����i�"y@���C��
�Y�*�A�y˱�0 �;�y/��۩?q=Ḱ_�n���p�1�
C��ۊ?^_�G�
*1�0:^�@�$�C�D-ڞЅZ�A���D)�nˇ����j>=���	�ULN����	��x��U��H�����iֺ�@�2�;��1���г�m�C��U�;¼�_b���l{N'��x+M�#�Dn��B�yds�amN���t/*Ǟj>��7�	S����a /fgTrj��ጼ[�:�7jת���� ���K�0fc.�_0�.P�X��xN��\$\~��a=��W5|$�v}�'�8DF ����qIE��?�/����ظ2�=Ϡe���ϣ2� *U���K�v��	�� c�Ѹ�(�k'� ��T�A
��e0#M�^��=�����Y�Z�6g��9�8�<h���(b���J���%�m�؄�rDQ�����Qy�5J(A�h ��[N����j��	��t-aD'õ���B�J/�oix?���X�:5d��7NfE��n<V%��<�������E�
(�O<)P$�--M��@����9��y>�NQl�l��7�c*u���e����D�jܜ�r����"���qbF݈�6$�]�!����A�e6�R��h*�~Y>����uxV_����gZ�5|/���-V`��go����7��N���<A�><5��iQ�A��ɡ���85z�P��Y��4�K2��M^N��dQ�eK5j��GV��A9ҷ�6��*��1]��Њ��5Nk_���
*x��,��L"F[jʊk�2��b��T'c�N���h�^��F�\i�A=��cC"S;K�oߗ���-LL�tAQ;�ZY��M�$��۬x�x&#� ��QŢ��H��Gvʨ�GT���oȈ�*H�7�`9��q���4M�|)	!9㹮i�V~	��,Yq;��}�O��ƈ��٨���
���L
Vf߸���u����q��i�|ƈ��Ʊ� ���e�#Zz쩕��er���F=湙WP*&����Ѻ���� 
�
���1z	i5�(O��h����Fa��;�}%�Di|���6�R�5��|��۸��P���ߪ�EO���
k��U*���>��9�" �����wű��6-�.�!Vi�~
�hǳܸ=OMO�³SvI\ƗrN��W��
f�=]38ZK��w�8�nσaQ�uַ�+}x\|�(Q���+����E�J_h��3��k�NI�[�<á����Ώ�%_����t��.5tw>|�����E�N��(۷���̵	t��c�F��n��%� ���<�����=>��)�����^/�=��d�V9��x�J�Շ�B_�m�e��K�olKnY+}B��ݭ��`*��V�������_jBn�j
ۣnm��{W��\���RP��ܚ֥���jU�:n�ZAH��ZV�|�$.�5��ͫl�x���5����RGfZ��qNq�K34HX�!1�uN�v
rto��[�f�?8�0�׮�
 n�|16"�o�
�B)����W���׫��V�!�K �R΄G�E�G8����w���2�O#iY�'�%p��}L@W�� `W!s��f��$�����V^�2Z>������+S�RJS$���(=j���p��T�lUMm���{��*(J�4,RD*���G���G�wd3J>(��K�i� =����%���KP�i�߼��eg=cmҹ��O��}<F7����* G�XUwJr���@>���=�����FA2��ϒ��Oӳ��ѹȭ���J������`�(��<g0��|�<�j)竎:����,�LB���L�K�}a�P5 i�"�Aϩm+��jWN�g/����kD@bGe��?�|���zZ���c�u��焭��7��t^���^�}:�'��ӱ	����ޔյl��=�ye�t��dW	N~Lf'Iy�#h��y=-�\�CR�bs~9�y�l���)Д���%�f�w���h�ħ�g��|H��.�p�X�>B��0���H���Yf�Y��X�U�pn�|iN��XS����B��5��Z,p0vk��O�P��F� ��%� ���ь�Z�ɕs�ΐ�����jض�4h);���A碷Z�":���|�uCt�D�D.�����w��l�Uj�Op�L����������H�?
*��"�à�e�~~��{l(}G�Pm�p�<���k�쾰�H] �\#i�ޛNvR�V�Y��q�0�˔���J�45:(�JYϐ�qA��D&��ԹOA0>+s������m_�?�ՙ��'�8cA�o�b΄��VF'E�{���n �RU>n	���cTF��)��ak�N��SؾC�[�ʪ���re�2�T�Mo �� ���	gN��7��υv�%�H;�&�'G�xC�n���~�Z�M�](Ǡ���r�RjD�d�z��Y���?��F;{�w)-�j����^:���i<�<����5��ѹ���W�*���"�+�GIo$L>��`�ذ���7�o.��WlE��c?W�f~Ub{�s�od�šz�M��W<��È���JCT�}����Q�+򁏼�
�	T��ei���[��4 �೯�>�ڗ����*e�v����}o��4������]���\����+s���9�I��� ,�C�(�@�&�EɂO��\��\#Jb~BgR^6w9����/7I�eq,t�kI�����5�D�{JT���s�a�h�F��9"�Ixy��4Ꞁ1���\��n����#wK����4s"��[������{��;�[h�s����ҏ��Č�nO'X�U0_ ��瓑w�CI�����N�ą�@����y.�K���o8�a��f�okf�ҭGL՘�9?�WgX���]*-~m.�.��d���<I�f.X>�;��u�P̹Oه@��78`�b�P�.����AH��0��������C�+��v	+��'�^z�\a�1���Gl9��. 3x�Ƞ�E�� d�뜑�'�&��A��u�XS�v���6TRU>��t��,��$�\�P�{��l����_tE:ڇ��w�-ݾ»txշ�6����j�.���QS6����U�y��ߔ�yH��l�������C@q&	�pi������J�X�>DV����g��;�?0�ԏb���s��0TU��1�.�(��y@��ap�A���u�/�4p2Ma� %��;$yf�R�&����'�%&�ڈ��#������8�(A�	���!R|��ݢ�`?���QYl�I�8��E��G�2���?h���P�!��Bg �`'>øw9��c�N�I��e!H-\/�hR�Ǎ�`�-��~;UMd�C���A��ߠ���H�U�� _���1��¬�o{���-�iI+t.���k�Uc��*z�M��������I~�r�4����qu�-+�g�N���(4-���l��1���^�?+���3$E-}���E���*���T.�6
\��[8.�9_�*�Ӛ���d���Gl5��F�f(���ۼ�d"��N4�wVB��՚�d�J���~��O�L�*A=P�6�+eɰ|~���Ŵ��������y�&L�u>��AVS�zA�`�Vݤ�Z����i�����pl��mv=f �M5ht/���o$ڝ6�OTM>,Z(~	�ZV��H�B������Y�"jW�ہ~�93q��BW�v3�@�$`[���� ٕSd��O,G*�h ��Zsk���㜏�R��>�j�5�`kd���e���M�Nt.�x�^yRYv[�r���AS�m<�Hk��'�-���j�I��ԍ8���}�.���ӱ+�������{�����j��0�J��l�A{��S8�5�ǊO���r��e�z��>㌟��&��x�4������c��+]|��p�o!�޽���茶է�k��yW+}[E�r�SdWO�R$�I�s�Wu���Z��F�J5��:���	�<��H�܎�g(h��[�1��ZgQG�V���P�>�z6��4t{�h��(4N<hf�ĥ]_�	*�Q0-�}|�e�vJ�Y��Z�VS�rԢ�w�-��!��_}�{���RA���7w��������/�W��g��%F�2�n���f,u��V"�)&�@��J̟$���R��b�uT�d������B�������5��sI؏�����>�����?�Ӊ9X��$�ɠ�&��:�Nx���.Z��8ڊ�e�B�u�G�v����;G�� �)=l�T��c�.a�5~\�� 
���Cw�y��?�VK*���k� �Z��ڦ7_��{�l�ᆲ�1�[��&P�(\$+��Z�6g^Տ�YKܿN %g�����Bps:&���V3kdw�g.M`s���5�,bAlO�Bҗ�>o����!�-��S���=�:�$}.�b�
����¯$�Yx����)�ߏ�r\"�P	k����_���vL^�NF�zFͼ�A�J�ӹ�M�qY7r���'��.l�M��DQ�J�h�
�5˾�Ee3��3������G��,�)��kkԅ� �t&(CCJy�e���e�a�KmB�g��3�"�ڧ��s�"s��o 5k�����}K�=>��Z�Ǝz��f�9��HÄ�S�ü�/���3|��
��V�ߘ���Ci�/tX�:�]�����h� qaWhV4�%���}�$����l�\�<(�2�͍��oJ;g#+"yN���s�'��S{s虻R���mN�:�x��5߁�(��ged:�i.��k����⨮U�'
~u��粿�u�\5�������*l�E��Mo�G�mg��d���Jؑ���l櫅��%�ŏ�hqd�I�u���E�-�A��vy�s<�o�'Vf�wT�h�;&u2���^�ɩ���F�ӊ�z��ү~�G�gD=?�N��[^v^>Y�(彽&|-�n��r�rݞ��i:Q?
2d��sY���6 ױ�#4�k-_����R�[GMb�I�bcF����*�WXE��Q���+��c3�vQ��}C�J�?�*��pA�YZ}Zj3��I��]�ժ6L�2��7tze*qv����KO�GOp���NcZ�
�r2_�h?m&AYg�CS�F�CB=]c�H�]�#H�˒l�Q�b�
���_�3��mch#�[/����q�e���;�����C�t���C�$��3��`��p�v�E�97��z��e>\\��d؆�������i���l/�����P$����#�ct�7Q��81̲����<O�I=XE���`5�װ�M��.�� e'Q K���$�ܿ��@��N���!�hG�H�d��~�饺�������EZGu�����Eeqv�"2��3���VG���U"jm�#"{�8�W�>�h�J�F���f4��n�M��H.�/XkS����EFJ�3�O5��WCr=�\��8ᄮ#�q��z�Mc�>(�[ѕ���&�jt�5>`Z`U�dZ$2�l�q�cjn�� �le�N{�L������H?�ˣȪ �)7(�-\='޸ڪ~��a��N����F��KMZ�ϔ�oa�Е���B�J�n��w
gF`�&�X�w�� �yTy"=_��D2�B�u+��,�)�Jg��c*:����s_�s苯�9Sq���wQ$��������Eth�R$�̘[Vx�Bğ�r�ϒbǉL�1(.������t�r��b���Q�q���Ψ�o��S�Z^C�u���ǣS�L68�3�R�UUk���*װTt<7� 4�ѽa��D=T�ls�3@��~t��J�I��ц�.���=��[5QjA�ls��@R���Kx=��ֵ�6��gK��VB��e�Xq"����=G��J/L�L���m���,N�\}�{*ǘz�g��h�t����<��H RS5ڦ�J�����|	��]�� 	֐_"?o��0E��{�]�A�P�Q�\���\Hj����E���8���O���9��ν|�4|6!����o�k	x�"�	!l�yv���b�3
��'��j�5I�/���u&<�+I�%m\E�!��5��$�t��kn�ͥ���q���[���d�I�� #$c�'�#�lvy��#�^+5)���Y��:��y��\�>v��n$9թp��=�;��֖���(:Q�6+�T�%�:��[X�����X�J��0�S��Ne�Š9�Q	 ctFM�V�V���*���@�SpYG�'ֺ�oD�:S��ĵ�넲���k0�p��)��%v7��%�M�w�D����#/����9�� �7d���[���	�^>_UuކkO�:�nu�G��c�}�m�W]I��A?ƽ�pU�V�x5��Ks���;������+�!�+�ғ��4���V�̵tDb�e\�`���L^��Ő�W:ۏ��,+����B�*U�^&75Ӹ���S����`�R�֧?����݊��mUl��/�����w4�F�8 ��0_�/��O�m����;s1��^@�	��A6�S ���r��a� �=Y�U�GF};߻R�*Rw5�����E �[�D�M���,�Ew�@'��H��{�U���M�f=y��~�3��c���x]2i��zp��;'�2�M��8��V6+�\���<��	�^K��Wq����Ӷ��Z�����2{��l���5c��B�l&�?���ՊWf�
�ڄ�ݝ(U�0���&�#�bb��5�T�LL�o7Y5@�4�0�ِ6U
�'w��6p0�T���迤�u�צ��j�\3����Ǩh��vEH:��+�Qtm�V�&�k��� 6�9�`,X�(����l�W����9K�v4��tp����oĬ��Z�L�d,~��l�BE�u��\�9��%���)�8vT��t������*��LMHe��R
���)�j_��f?�����|j�����X���y̘��8p���U��S2��B5Y��%?�o!��y�M�_���Be�4v���û�{j���4H.ߒ`a0 m�K�ˁ�=��: �nַdO�c�Q���^����`n���u�o�Mp@�ŕs~&-?1�����
�PU7s~,i�9�9	Hg�>gD�34�e�GZ��P렖�%	���~
�|P�r*pƛ�@͜/\�`�7��9׊� O~�{~έ$k�`������T�V/I�a�����9���tgVLn�MԒ��"e3����.�K8�Í٪�|?�SZ1�iTF�M���!��bf.��7w-20�ʵR�L������渿'Cؘ���D%�,C��9�_&�/�>}������k��n.�l��z�x�W�vm���6�&�8�9����85ݾ0-�hzw��E�u5�|C�bضh���KN;��"�
{�@+��n�_R�u�s<�q
aK���BL�[�!������R?��B۲����r��R��jfiF��8����%��a��P��`f�y��+������:f�"ҁg��=N�T�������G꾢��A�ʳ4�l�9��k���I)��+,��'�4��!<1�x�:ϳ�a��#�==�5��5䤍���$�V�%y��n�[���`�H)ÿF<]A,�KȊ�/��� $V�T=��7p�RKѥ~�.���R�3�n<%�X�2K�´W�Q��g��r;�mi�I3�sV��J�KU�����_���-дmq܍9m:���P%��2S��46ɾ�=�k�{���4����0��J����7��9!.0n�~�a����`�4�{�?сhZ���n��?\'�b��=r�82���X��$iIC��F���@�X[X�;�����E�����|��E��Ρ���]㾔t4d�+�6��3��<�!\��y� H��Sc.(��t�\�Qr�wá�=���H��~v�Zy uܡ���g��6�w_x�󬸊�w�~���-B'��(�9ɴC.�kY	M�ȕ�����0i򷿖a�4-�x'���}�e��A�Dei��xK�}�>���M���e!T�ܗt-�����&>��߼p9�K��rh+'wJ��l橍҆���`[�me�B	�`����x�t�9G22}Ir(��	X��\w�Q�2~
o�Q�]~���d{�fe`+az�rW�zw4�<
C�9���7r�m�a-�;bNz9@����ȑ�-r^�\���������N�U����W�����"]�;٩=��t鄨r�^�O���m�� �<�eP��c����;�T3�aL@�<�*�4}dC�	�oŻ�إ���rh'�b�цS\\|D��!��1h�K7n �� O�RT�� �Qm���(Ѷ/� D6[/$,,��rv��l�Kc	Y��r�7Ԃ=���2��[Ϭͱ�gq�`
���2���#D��T�e�f�Vn�6a��K��n���R�Z��N�h�����)ͣ"��c��u��䨌,g����6˳�!ʈLE��y-��w@̉S�L&�=<�[�L/��L���xߐ�u���ɪu�bܶo3<O�C
0�V�%+��\:�+���!�)��܃ �&��Gm����k-f{vK1N|�Sp�	e����+M��r7M�6�Y*&يt��5/�/
�ߔu��N��5�e{t��L�	0����}��HX��*�8-Wɘ��t=x�ڹ$�~�FH=� ���p����M-q��/aĶ��ן�$
)qY'Τ�� ���fi#ڡ��B�ɍ�>o0�<�����G�v�K��C<v�����Д����	Z�:�Э�m��3y���۸��Qf�r �y�A�Mh.5ؑB3�ʝ*��ddIE��T�t��qA�R@�o� �TS��	uɎ������~�'�:�ﺤk��q�M�~� �أ���x�9<} 0%.����rb�D������6��^��s�~�J���$p$���åH�	��� j��j6Sk����j}^��xIa�(NÂs뺉_�UtS"@�N̠���j�ۢ��p�rL��y������3�R�u�I��.�lj�ԲL=p H/k���fSa{ҹf�(��r���Y۹e�=ę�筿B�󐇻!��?�q �k�T%����lIW$�qK����3ܵ��Od���g�
c�����f���+�W�R0�;��T��J��lʛ�z�x]�di*)��[�Ӟ�.�r�~\JI�:pf�(�ђ-��������D_P�di1�2ٿ�w�
�c��U��	̭T��a[�IS��@�?����a�A��6��eߑ����i�Dۉ�o��L��<�ҷp��7
kz>�'���nO�]�i��.b����Uj\U�;����
�c!�C'�*�'�=�~���u ��]���â���J�qk��a���B>$�S+*9����>NY������I�,���(@RȄ��a7>�� �o7j#�0���m�uŝ����G���$ѫ�Rq�-�r]�OC���ZKS�c����`�|m�RC}�ЮPr�S�zjJ������<���d�YoC�@}�F��ON�("��w)�#��ͪ8j|��H*�E�:��������
gu�q&�M�p<«��"W&҅�b %��L!+���V�4$���>g�/c��p�����rk�߀k3���?׺σo�i)9�Ӏ� Dlp'%�
0�_s2�~2+��@IPD04X�ؕ	5�E:E�B �w� Dw���V��߿��WČܭA� �}����b��̤�//�x7�g�ygbTv�`Uk}�UQړUʡ��m���772�~"��l��JΞZul��hH�����x�)B�ҌR6ECOĐ�0�Bp��7�eU�L�_w<� o��S0��JEtz=.�X7�Do�ihC�p��A}�pA�ҍ�/��>ސ���A(�� ���M�+��Ad�ۋ/.](�����
��%��f:l����ljK�?�s�ߍ��ص��Nۆ�\����m,�x�NkB^�����,ϲ9oy�T]+B����L��Ѐ◤09�FF��5Q�O�[�� *��P�;���Q��wR	�7�BQ@{ȁ���a�=�d�
�ޚ ɐt�x�
9�����V��Z�-�G�̱|��3/��/�o�]90�7�M���C��K{�9�zZ��*Ӵ�຦��l�R�ߪ��:����w�Iw�߷��}��\M�q? "��]툍ex�;Ք�.�l�K���J���6�8��T�"ImV��YE��]?���T{�3��N�`�w7#�K͵�.�>��eu�cir�Z�o��TO�3�1�]}��Y����!C���A}7'��8=z�O	+�Z ��+Q�U�Up@�Ѥ��r����Z�o��ϝcW�^ke��Qu�c`�ʒ�d��Ն�nT8(�a�e�n�\UY]���ʏ࣎M�9��Ϋ�
w��6�9:�ӟ������!gQ9��R����
j�73�������A��Р��Ł�#�L��Io�Z�mVB��gA�T�U�}��k�$O�+��͔���B{H7��a��+���ia���h���1����g�;N�u��t":�CV���Bހo�l�� �zIt�p�S��Ό�4�L��Z�o^p�"(���&yJ"��r�S�=a6�5�!��"�h-���ɛ�to�H&��ЖJ����|Fh�����7�Y��C��
�M�R�Wx�֪^}08gH��pO�+�%P$�J)�n���a[v+��� �#�[H��4v4�H����7�ZH��+9��X����㗫I�Kd<A�L��;[��}:�6�謩�=�F�Sܝ�ï(�P�_.���ψ���[��8m �8��tl���*��1.=�H�(N�J��ZQ�a>�f�5X��n0-�(=}4}]��L#<"��d�nw8���O.�[Y�ǱM��\5�N'�ɐ\0�]��UW(2��J3q���#��:%m����-�� ��eI|v'��hϣ�jN�wh�TRu���Zm��+oD�B��,��6���R&���($㬀X���2��!��]Z�����`�'����H���Y�4�Aj��cm?�B��v���n����.���'L�f!܄`���Z�G&�$�(1ת�/��.H��8����V��M�'xfX'�'n)��X���>΂��r�D�g��p>vG�J���I9���[���]���؂+K��]�Yу�X�-��\>�+����w
�'���>{��[�6�{ҁ�1����f�f����s`u�/t�?Έ:b����~����A��Y�~(�T_�C�(����>��y��d����
S���	ηth�D��8Q�%eCܙ٦) �e���q���,飍�qO�Ȁ�ݔ rL簕��>1�gBlRm�@OQ�W�Ͻ���X�F�* ��ߑe�-�o���Dk�][#���FR���Ｘp�8���@0�.�-�ji���Q�:�Z���B{W;�?m�p��d��r�b�A��*Xf�K얣�L�S�[�4�����VYM�V�����ꨨ���3W"���)��~���ySr��9J^xl0#���x+ޚ\��e&�N�Q������
�E2���/�����uϵ�^�����o�L>s�`�X�A�e�T��̱4�=O~�Jr�9�E�O
�G�.�����T�&-�v�tp<��;����� 8��lg��W�NR�M��4e��P��P�fG�,�Q�B�Y-C$�"�TGS �A�+0�:@�`&j��Cг��tFV��,M�H7vJ_3����G�h8bA�8��|^��r�NH��r��O�$e���>B(?U�`V'�Ã��	�>�Y2��ƠO�a&�L!��K�]o&.'e�����������f�ÂBb{�ǜm!��!��I�T�`�LvL����Tz!>*�eF3]l)�,pg�Q�T�(����Nң ��6���}M藹���d�$oJL��#�k�#~�հ7���1�yo���*�=az�460�+�w������h^��Z5�G���X��\����C]m4ࣰ�'���j5&�"|U���ٶ�3���O屻�s�i!\�z4����ڏ-$�.�T0�.`�NnLS8s xˇ���G���8�ku����f�`Er��|}�늲�����T��빍(��	�/y����·_��][������w- �;�Dn��iI$>[�4I�Ю�D��{�5��a�Q�},6�<�+ků�niF�;#]T;�$A�00��":�[��e`��_Z�iSu��G�
,ҩu.���C�#����L�K��\�61��������� W�[�6��SA�U@�+���	����÷����e�iGGv��b	�j�]YM���n1�8�icen�[����Oý״Շ7?�Xoa ����,}ƃ�N��,��)���ʘ�'�m9�Q��raS�uneMl(b4#�CuN���21?����ö̀>Q�v:����S�)�q4I�	g��!{x;��P���чt��y��c�:���"ژR=`���T�6�?e��碵��-j�j`I�&M�-d?8T[���8��%�[�U�"~�AO�u���ѩvF{%3�,6��ԑl;�L�hg�����R�W��-z�q���f8
Ѓ�eX�M?t:;̽(��	�%
nK�򙰂��0f�]�~[�����-�BSDw���rP �@������uN�1R�������b/cO��� ��~�R��"J$im&B����z��4��������2Bpv������ ǫ��%�*in[�9����M6e��՝�P�r^��VKK^9}�������!�s�0u���F�f�� ��E��)Ã�\[w��#Xn^MC��=[&�U|��{r\J_1iK`B�t*���[!�2f�l%�%��Hn�m������B��}�A��HkNJ�~-���_�y��{���3���Q(���]�`~]ꙍn� �=�������[h�C�He2s��ҥ+�]r���� ܦ%Y�Kl�{��4ȜJ��N8QU�����t�����`�lTӧ�UGQ�'d���Lr�^^��.]ЀP���}�����1�Yý�{��]�U�tV�o!m��Gt����ShM���n�I����hA	Fyփ����*��P�kon�O�Q����%�<�j���Jح-&�/Γ3�kl���,ɀ�>�������X��N��#���/��V���(z��<�4����,�ь�J5tcG+ŕd:��E���]�\9��;�vɀ�W��q���� �����T.q0(-	���
Y-u��>��5��-Y`���3aWe����MX��&����F(j4�[��FPAr��"^40�A�*��zJV��*�b���F	�}���J��R3mM���C�0��ަ_��/^���4:K vi?�'N��;o ��?[��k��5S��W�FlD����/d_Gg��17���mi=ތ�ئ->�ޝvW��a��f<OX1}�[fȐ} �'�G�2g����A�Kv�Q޽W|\�'�n�wp<�-^��ߴ���E��9��`)��HǼP�`���M�VNa���i,EKDP
���)0��J�'Tt��j�բ'q�-�S���][��g%l�N�?v�M�|��v�lڛVRQS��[��.����	B~I�7z9��e3}̿��kZ�|�L�s: p��>�]����+	��	��J��0�R�<D��<��j���9�F�����`?�4��{?�|���O�<�O��?�0�\�g�|�������Y�]������#Ga����*�1�+��feQ���};�}����Lxk�ј�v|߰pcf�9 AMO�<&:#���H�3�lPF��4"���!>��`��+�ve�;�����ef�&s?n�o�@�� ����K�^B�=�H?� ����5>��S��Ln���[?\׌��Υ��W۹R\�~n˧O���CY�|]�����L�H�,<�5�
1-��c7H���-m�3��Au}oZōc��� �|2�G,��*ʦ����<ǵbp�����{�������S�A����`]��Pn_��?�N,�[�)Vd<�S�*x����IY�p>R��K)�����ü^�09(�|�q�Ɣ-:����BIF��O�v�4��n�Q?��`����T�dͼ �Ak�<����KS�O�G[3:,J�yl3�cg�a��e�9N�(���"��Z&wr�-��bJ�;�'�V(��G��pk�:�|rZ뇋�s��=h���O�
Q1P�Q�ώn�V�Z�|�_�6Һヱ��.�����ե7ck��E�E;6^"���P�\]�`�����`��b��N��Ý$��k'��XҢ,N'jb/'�ۀ_��\j�Gu��y-f��5����
�"j��Y.'&�]|�L
���<�'�E6-�-I�%*m�eoo�͠���A�&�t���P1�Rk�\�	[�]�2�܅�Y�L��Q��2d�a0i������I����[����څ�:������<�ץA68ԫ�_����L?�XN��E@]!�'l,�����sLXF�uQV9����xm�3���W4x�{"�n1���})�Dq��CM�SJ�
#I��b=�B8��C�F�ϗ8i�Yu�oг���,a΄i�X~�]�+QC���T��h�\qNa����:% ���薧^��ZхANEU\��VWs��ih�.hiH�S����w���3?��K����hEc)��0�+v�	Ϳ���DK;u����4]���l�[�?�َe?Om�k����V0Oe��\TF�珍�Y�$��$ڥ@z��m'�˯4�s���D_�Xl�ON�AC�42_�cE#�/�l]s�u¡�ka��S�Qn�-ժɉ^퉏RU��U�wc�h�ŕ�oHq{��v0"� $���az[�K������\	8���P�Hb��ML�DE*�'_td^d��̈ ��4ɫ�6c<���� ��ҫ[�!���y�Tm���닍�a�{�q85�;���z��8<��Q �Z�RBK�;�MNK����iU;�FM�!��-���� ���Ēr�[�� 6?ƅ8��+�JC��=���)�B��棼+�T��X@u�羠leXA�f��KNR��PK��:��y��]��'2MW'�~Z�}݁��bWs�K#��ÔO���j�a�w:A�lMC"�-�#p�)���t��D:���+� ��	W��U���#��/��d�Ն4�$UI뾽�tJ�;�P��WsV���L4cxé.I��vv��&E�������f�����B.Vk��sHW������S����߈,�+�f���E��e�E� �+�{}���J]����,G֤��u�ɜ׍�*w�F$O�P��O��!Σ_��Z�e֓���N�fޞ9�����啉^wsy#q�Y_P)_1.8�h��6M���������8	KS� !
FD�i��Y񓗎T�}��FjcP0��`�55��M�ȶ����G�VM���J�L4�X���3ez8t�������A9���1���;Y��Nj9�G̖	\E�}�ӑ'��d���ok��gO{N��~����9ՇJ>���6¸�W���e����U(v�rpܓ4�6L<=�ӽ�?�|���fj��}�n��ȍ�ENZ�Q�a���a��*��x����<YKB�O��L�~&m�O���s���(��޸�1b����Dބ�|��SC��F�A'G�%��5Ｍ,�A4�*,UY<�w�3��
������	c�\V-9��P�j`�+@�����4�_+J!9���YfR�e�乫Ǒ�~�E<]�e�
���bo`Q~�@�����Wܯ^b��פo�]�9�G��"|�*K��sw�w�R�>1�"�(���h�n8<:=�`��g�K"��u�����+�]?Ƃ}|;<�P%@�T3�T�!Ԃ^k$��`Y=Ip&3y.��4�Se�:��$�!(k���ׇ�.�;>�ma�5/��'�dk|�e�_.W�Mo�^ܻZ�bz��:�!�1t����U�1������%0��1]m��6�x���6½��n(Ǐ5�f�I��,FtH��[��mI2�B{�K��e��׼$'B�92nUjѨ������@޸i#�h��M��=��ꋪ�+�a4h|�-(�w�!��
A7y�_b	q�fw�h��-�#�|(��+�}���H����*��%!�\�{K{Mo�4.�C�����Rk`TZ41�kDq-~�|���0��1��p�=��e���q�)DØ	�|�0t]���^����ɬkwI����x ���3��mb��a��:��9��[R����4����u��>�
� �	Of��ze0<yS���Hc9jQbD��a��x�Q	�����w�*���˄ա��֒���8���OV����ޗ!��5-�w��d�_?��j��yZ
��a_��+G�N�詑�&C�p_�!��R8N�!���<���O3�~,��-�
KV��=f8�W��Ff}�O�B\ī��SjV�6��ט����	�|IGsZ`o�BQ��z����a��{�,rW0QX�����)����x�(-���3U��Ze=�'M!��"�i%K�ҌS\]wuˁ��ȁ�r2�����mTf�l?���R\�:�k�%G�\FzJK*��-Y�u� ��~g���7S�:&��U�,|�� ��%��������9L�Y5���KDA�g�����A_�L5fL�x�T��ͦ�9�/�����s�<�z���\P��r
+A�C�d�g��XD��x��M���*�tk�dtİd�� /��-!߻q#���CN�g��J3A��Pn�"+UX�M����@�&8[�m��2���Hj3݅(D�"����)nǋ���WCDc9H��sͲ�
�4k���J�*oJiNkBku5.�O5G6�K�VE �z���ӫK�*���%��8��A� �����LXe$h�mKkb!���v!��Q_�x����Z��M��s%��2t�}�7M�έ����)]��=��;ui���?�<��Ϫ�|���=x���4&ʽ�d��bo��if�pBVh�{�P8w��/�mVH#3Ϸr�G
��nfc���UCn�x����S��V�J�@��;�ʨ�����v$oG�N�q�Y�䭂ۀ�=��q�z���p݇uu��A>�_����A��(&ʡ��%ډ1�}�*������L������P�~7G���֮lʖ���ڛK2�dӁ>�%'l�l/�.��$V(��7MYm��e�_��%�;b���57^���-�L;�+����[*�n	A�%����!̺܇�l���{[l��gG��4D���K�7�����(ȬW[���A��;�;���1�t�M}�u�׫����^dY�o��Ng��#҆[��y/=jJ�}6���4�!1+�ϴ�x�w��� PD�}O_s%��� C&j��y����~�o���k#��-��C��+�s���Oj���k���������񽧸��6Y�9�:�t6���K}�����o;��=
��H�{_^�;W��|y��ł�S���>:���_A2�2cS�f`��Pפ����i?ڮe�Ų3FX��?ᣜ���0FI�"��!XC ���\��:|+3j�Q+�0��?$���W�	�x�����D���cj�Q*n?+��1��0'�����p��Y5U�`tQ,z1����ԟ�,��q�2""� }��EPxĠ��;�`Xb�@�q����xF\_oUEajj^��C�ށ�|�s�#p�2����dA��� s�i痒NȨ��|����'����d,T�G�[�� ��u-Fe�S��s�ħ�n(� ̩Ⱥތ(�A��3Y��*�?�������#ޞ�M*��������6�a���k�Zͱ�1�xx֧�=ww����le��s���ԓh�(/G�������>
f-�L&wI:�����!v���=+�=��M͢�0 rX �~v���>[�)��\��p�b��:TBM_n;�Auҭ���lo��j�6e���ڹ�E���H��\�:�Y��fؕL�N��MH��#���n�'�T���0��Yx��zv��z��RЃ�{	����`�U)��D�e8)0'd-M�i�2L��"D/���n+gt�SCGw ��R��t'�eD;hd���Ӽ�Ao��o���|Q�nVt�(�i�p���_]Jhh,8@��]v�����қ�=�U�20f]���K _�kh�f@�[�(����W5���t��`���?؇`p����9���d��cޔ��(�hdH'.�EH�c���G�՛�����x��_q,vgN��K�qfł�d�F�����"YV=ҪT�쾡���(Soj-�3�����cB�8��9�[��w��BI[/���K�n�P&��L󹤱���hJ�K̮ă�MzF[^0��1���������y��HF}�K���J��,r�\o��I������\Y#�V�^8��� I;����+�mMR&4`����(��n�U4��N�_�����$�Ү�Oǔ2�(.��~� ��S����S�/�sN�~��C��B�TB�P{��C!{��X)�^װ�U���U?�1�.�|a�_ǆk��a���y� ��10�G�9�6�W)�2_Ucn2�wM���׊S ���Z�mnE��">�⤮k���H��WD$�CFaxN3^FLB�;b����᭼������Hz�%=���%B<(lǃa�]�l�FM�Jx�H�0�����-��cXa�������"�K�QT߱+3�߾��q�|����?z+�6:��}~b�M�/�c ��-f��W�=���i�1�)@D��I$�Z=X�~��έ)����
��z�i��4L5�ȝe�j�J�S�G��fw�廷m���`�f\�>�h��.*��>`�2���4Y�2[g�Q�>"�ƛ�"�	l������n�4�!�<AQHȆ�5�y�sˌ=ma�����[˖A���%�(���D��J ���?�\�(G�IJj�+9d���9`�Pύ��ā�IģM&̺�D&t�ݹ��z�fJE�L$��9k�x������n 9څ�P?���LLZ�⫮�I����3I>;ppu�bF��?��v^����������FHa����"��8L`�sSe��,E��b6S�f7ih*�$��B�]��әS�\�_�.a�q����������#�Bn�����m~k��~練���o]��g���lV6�М��\�e¢;"6#�G�Jx-�O�buhg���	H{�|�DbW�lZ�7�i������E%�Y�\����Gn�j�4�Kh:�
�O�!/�����7I�!��=:��p�����r�kӏlp�EÝ��~�ӌ�;�[��OZS�I�1Nľ�́��0`Wo���3���ߑ3+(1S�Փ-߆����8#Pu�5�$���f�.��n&�F�J���#�X�ҷ 9�C}/�%�@&}��T������u�}�ͷ|���LPo���?)ڙ����T)l0FV�w�e��n���(+�����~bd"�����9�>yg��&�a���q�w�0��C13b(��+ɏ�%q�1�<([N��i�9�����3��H�"%=���8	���9��}O8���b��V��6��w��C��i7pԜ-]�)�՛��2���(�kf��=�l��T���'	b����?e���ٳ`�ф��j�rR����n�T����R���Bv^���	��FEe1��39�X+�������Щ�Z��x +�pL��Ǵ"?@4���P�CRP3+^��(�!���i��M�o�[�-��L|�P����,� ���KJ��8����J��ri�{Ͳú.Qu���N ��+�$�#\J:��n|�e)�Se�?�?M����+�Y��JS�v%�gY_Ǫw3�Ym~�9�|,�2x�:�N-	�U��m��7�D� ��^M
��[ž��;ʂAS�%�״z�^o�ҩD�D�J�N�����(������u�/��W��sØ�3�����:��)�@�t�/�c��	���d��?�d@�͆Q�1"�[��Fm� ���Og�zZQ�����͏��z����W���w�&�ױS�o�yY����Ը����P�̧���懞���CY�s�*�R��]���fq��C,�Q���*����-E�����r��h�������%=�4�)��eZgP��j���-�_As�Y��G� :GEz8C���$e�*0J�����a�T\���l!��2�UV�&�'�v��>0Б%�0E��g���%VN,׊�E9�۷��:Q��ʴ6R���Bz�|�����+M�����p��������� }�l��;���ń+B����R�a���Z�bMNo��o銊��:�!�G|?���,���
R!����ky<�����Y���dO�M^U�w&e�����Z]�clϦ�� 9q���t��&9�KT:��[%f��I�z��k��s��ʸ(�����;��H|!�CM�h�?�xh�+����;�|������gȿ8��d�F���G�eP�����,���F�Oޢ�F'����Z���J�֫�O+'�����ÖY�VD��B����n� �k�U�P������@�o�_�=P>p�sZ.~���Y��6uyV)�m����Bb���۲j��	'?��9��3-�UWaV��W�ch��[\E2oD�
n������`��be59,�8����b|1���C�CL7�x�i�.���Yr.�2��<}H�9*����h��EC�_Gglv.�i2�ұ0�r� ^/+h�����S,I���o@���Z��僜�$���8-��<H�S�"���<�rU7f�F�p_>�u�E
k<=�J<"�A۽���-/��'�K������}���R��sa;��?3$J��o���h}�<���%��*'GF��i�nr�Ry�&n���t ��G�m�1��xi7R�� �.&g"~i�m5{F۰ ���O�
M�I�;
*D%��4;���3V�%�v+��?_�v�)
���`q�L���^m�s*�J�o��y {��:�1!��*����tjO���8��/�6�GѼG9�4�ۧp���i�O�Û�j��X�����h�tS>�����^���#�'&u�s��~fq�sϯ���T�ƣ��o��L��@�TI���c�f���W�
i��V{DK%�|�T�xX�?-�W���^����fD�D8M�K��F�~�����e�.x$���_2��`��2�3]o�ه�!�a��~J�D����t(�Xy|���nк	�"-��U�AC����)Z/R.&{X�>����Y�r��+q�5B�J\e�?"Ψ��w��$o��iC���ӏr���$t!��k9����Q�	h���!�O	��䚊8�{8N���&�-��0;Ͷ����o%�|w�{��: >4t������ɸr F2(���&��&��c^&y�	���4EΦ�w�;��t6��Y�S���1z����+5;����5��B�hz rl2=LzF?��n#�`�n��y)��p�K����Ggx�o������[]4��d�˰�2,҈����U�2kEb}x�/��m'�*�J_�������w�l��id_�����R?cx��
A�4��dL�+��
��U }���f�g�����ٞW�F^p��K�����FԌ!VI��hu�k�>��n�˥=9�v@Ħq�R�a��|?Z���H;	>���T���RE��\���d�Ll�1��
~�;}^��wz>A�ײ�P��|㔓���/|u?Z�[u�F��U�Q�Ն���ߟ8K��VJ�_�6�0%�C3w��V�1��
3��Um��A��`��XFE=!��h4�t��/��|�$�fT9c��R8(僮�( -���$壤"O5?jRWI2-�x���L��mtPd)xP�@�r���Z�#
U�Qx�t|��S����[S+�|�_8���¼����Z9���[E�Z�[�8w��@��fQɲ�=g�tI]��M1�.zkcp��8�4�]��ߨ��e�N^��k�cKFo�*{8F��]>��@�o��	i�ݪ�,ڵA�P�`[�,�Rh��PiC�
�oѫ�4�� ��s� ��P� X�Հh��嬈�=��_�0�6�Vh�B�A�}�;��eS����02WF1��e��[>GU�e�N�ŚG����t �-y���I�{���ѷbf[Zp#s�k�sNgC�Y���!�<�Έ{/���Q+Ħʌ[l����f�l��D��q{�' ]r^zXHQi����v,N"�JB�E�زX\�{��_I<Y|,垄��\wBTb奬J	���&mI�F�?yX�7�u����߳�"���;h�|1v��%�������(w�'�jƮIx]Ti�m������-0u�v�v�;�\q�\����,��f4zǜ{�ӥ�5>����� 8H����.�5����j��'*f�H��_=�s�Ŧen��U ��rK��2�4�v����ʝ1�ћB|�h�4�2paSMͩ/�K�2co :�Tlߑͦ��{+4���7�kC	�G�2����8,1��0������ ,�9l�e5R��$�뤹�jYs�y3|�a�����y7	�o~��8RE�}���b�v�o���Ѣ+��)s6V��N�v�E)��I�<#H+�$�^�ٯaEٮ-��V�ɂ�#XV�l��g��dܶ%E��R�Q����/7�^�����i&8~w n�I�bsiSog���0��\�I�D�|�g3nl�Oh����CN�R7��*�B��3�XtW_����5)J>b�k.��H�l�qy����J�sF���?�[�r���D0^�gN�,#;Kø��v�8\�^?��nۺl
��.
�����O�vk�
��Ư�|p�{m���"�����i��c�KL�	� �����i��0{.�ʧ@�R���TaW{�_:#��?�$)8a���HD|���N"-��Ekf�)����V�a�Xg�"8^P����}&k�r�B�?�,N��T����mԴ,�L�*�L����1�;��^��(v
��P*�+�k-��ib(�4#�V�.o�0D�~9�?���s؋�܇}K�:|�կxO�W�q2���'��A��^��۰��q���o�o�� WC$�A
��\s���N����!6Y�~o7���YG��%k�;�*�4�'��n�u����w���8}Oj>=����M�g�n��:���Ч:��s�6�W�'�I�^R��Zf��a����w_ _��<}���QQ5>g���=) �c���1Rݏ�IX�T+���7w��)5�f$`MJ^�$*@�=/%{5��δ>7G�U�aCy��j\!{�c6,��dN柫���Bc/�E����aI;��\�_���/�z���:\10�K;#�{7��1�,�O��k�b������|�'�I�-r���@Gs"x�iJ��EC�m��nG�.�lNW	?������=�!�P�}�/��@�:�-*��/Ȝ�Z�>NZ[�r� )��L��0'S�A��1�p���g�	�-M�Eo���+q�����O��U�	�A��$s@Ӗ�r ���ЈnX�D��E~έ���-������Γ��tQ6�n5��J��b��FM�a�4h�%],
2���H�����]��|O扢*��E`P�`U�K�?�J��WS[!��ӽT��Lu�l�S�.CyM#/5}��/{.X5{0�k%�JubٔV���S5�T�ص�����'�<���I�l((#b�m����a�l`AZKD�䉓1�PM GtXXeF*�k?����*�2�USww�Ɨ�#�tFK5+O	򒦤��C;�%��oA����?�������c4*������8�D������ޝ����#U��s[�Z�+��Ò̓N(������꛺CE�n���n�I �2��
�Y�}͜����}B��P��\��ɍ9ƇIDdK�Ǵ�-��f��l<��Iuq��KP��ޔ>tTy�E�o\�q�v�oÃ��i"p�Oeb�OSC��k1�o�|P�]�%LZƞ#D>ݢ�8�������B��>�;���8�q�f��s�O�-��'�cG��,�댫u��(���9X����g��7��}�!=�$� ;M�lZ�Yĭ`Rl.e�=���Ѓ�F�w,}C(�:jRԛ���4tK���hߠѫ�|�.�����c��4�E`������BvƊɢ[�p>(dC� �4�m�6;VX�1�g��r)?LC��]��z��L2��<�}DG����Ӂ����S�%���l�JU�ŭ����{'�@�ڥ�AK�t��
W,�͂�R��ص`��bw#�����F%I�t���?+�v�����86�A.�3=$�{cJ�Z%m�������ڕ���>�%d��5@�^aheS�Xh��Q��C/����J�~w���Gi1��.�������^>:�9P��N�>�Q�$[K���J�ܺz�le{����GE<Ʋu���k��N�����1I���ѩ����xݼ����n��2���̴Z��j�c����f�5�iK�Kx���˦ԭ�6���^�b+�/�;\T��i�tn1�e-co��:(�WO��s��T*��u�a�����b�t
�xJM�)�a���܏n`M0]�R���1e�jo��(�C3���8*69s��@c����n|8Ő�v/��N�O7�c�p�������Cƥp�&�6L%AA��e�i�inUib�K�Ե��$O���r�[vNӧ*J�,Ms��7�Fo9�
5���ნ�" n��g�T��t{y}d � :�YFg[M_T��{$��X
[�Ɛ��p�Ϭ�+�G��#!:jU�Kk¾�����i����6w�� ���Z���}�xg�b�Rse�2,~��-\���ػ�c6L<�x��Zv��c�����cÉ��L2��<$�̸�d�)�V��h*� ���l�@;l���~k79ͣ��M�U������ʥQ=�L�Ө���ظ5��p�|2��6��B����H�72^�ټ 	�n"茫AM���Ӆ<9#�5@�*_�k���2���։
����"�d�.k������W>�_&�Z�wۋA��^8r |P����W�D�)��/.hHRI�2 zǁr��]��7�f��UW������C����k~ 5P��p���������Ibbc0�䂌�g�'���(���"3��>����\�@-����P�9���*���ayj:l_������%�����\���]p-��&�re�+6
�3����8���g�!yy0K�u��Z�B�n#��򣐊�U�Tq+�Q:1�!�,)4�����%3m,)ﵑ��G��1E�\$t�, tȡ��"r�lX�&������^J����y�!>�F�ɠu�&,Y��pt2�l)F�Kl�%*S������Q�o˭�k$��5�IXX^�ɡ���P��Ϥ:ۨ�|txҢ|�q�N:�1i�`a����C_�s�`��ہ`Z�R��||	���u�&<m��T�~&e�Hh;Q��1	�7�E �&wϋ9�ޮ�YZ͍r���tk{}<9i3��K^��$ؤ����7	���z�y�J�!�s�!�t����_Q���N3k,~�%{Ui�)�#��>�kn6G2
�	?Bp��D{��e��qە�Mo�"�_�o7�@x�����U�9S�{as�k�80��a+E� -W�+�+kF7�pyӠ|k�.;sj��i����ar�NT/7��I�RK=����{�*�R:&`[���|{����Éev~F��<���z�K:�j������N�?���¨86��3MdEg��Pӛ眘$O��O=���*6�鈌���+�������PiS}jv`k���%�tnK)?KL��-���Y���E�����M$@���^^��	�^g�$>��%�L�R�"�`y_�o*L�z���:g�X�lsS/}��9�Z�g�0x!G#1���T�ǦϠ�)j��,�W���o��0l�T���	B�7斦i��i��g�K7b����T��}#�D�P��Mi��+4u���\k�d*��iT�����М��۳,7[�nOE���i���Ȃ�qY��C�T�� ֆ�vo��8�D�W�Ä=����f"� �TM��g'G���=�ֳk���E(z�SZ�b��N)5�_�u��2�]��b�{�-�)�Ȁ�����1�p��{��ش�����\�$K� r�ŵ2Z	Q+_� %��gj�6�i����1
PV��1�d���x"`��HI�X�����g�.]�q�QA|q�qi��\K�c����
�5�E��#�A^	�\kA��A5��`��P�I0�������:�ZO�o�żj�9����$=���nf*"�w�t�ޤw��519���y�ѽ^����:�o����x���3��&�+"n={Z�eq��Xc��c�s{�Ca���{���wo�@X~Y�/|�w��c{q��aj�Z������%)9N��'	��P2W�Ԡ �%���'�+������?y������N~����E� ��U���������hi�J�-u%E˼y���%����≚�"�:o�h_�:(��r�4kI�bt�;u�n�ZH�Z�ݞ�bS��;?$B{ȣ*V���؀��U2�)O`T��k$m"BK�'�xB�yJ�%[zx�P>z��Hr}:��iQ|�G�m�p��o��#�L�"�Ԃ�p�`!�����v���}97���ɧ|��<F��hl�d���7d[!���(BR#�;��9���7��O[���ul`.~%�}� `h�m��>#\G\ �T�<�e(uS�=��!��An.ԥl	��Y�n@�]�U~r�ݡ'�����Wʀ��۾0����W�݂���r]�v�YȮ��ǡ��>���JYu��]P�N+���s��\E�Yi\��`�O�Dw���*b-��`L��I��遴���%d�!�m�Ra*��톏�U۩�hm�.��7*���Γ��9f�t�}#�\��������#l�$���T�v�΅�i��'a��[���Xl��l��j�����sC}���9������lyt�LK�v�
�n�X9���T�ܞ��R�z�a)�::�L��^�d<��Ȥ��㣌*�s"�BZ\+Ok1�&�m>0hn,���|)��zӢ��&�[�8����w@�3�:*Ѝ�Z'b�ۓW�$���`�� �H���i�k�R���z
��b�^6���� �s�A��KЦ!�Db��710���C��50�Jh*���e��=��풞F\�̲c�@0�!T������"S�s]p��hN�.U6�Fd�cu���b��=�o����d�%�݀�������P���A��U��JOҾ�����S��)�ѽ��ApҬ$���$�\�t�A71���mwMw'��
�^����/$�ln'���R���S⻩U��b�x��d#�"��S���2��bfB-�t�X��ڮ%b�, �x4k�o�ȝdG^�"
6"Dap�
exI
ڰ\��f�e�o�2�����|c��F�[s��^Y�����ռ�C�,r����;��q<G!*�y �qby(AJ��/jk�����'?�:�՜��oɠ(QK|�#@c�$�
8�7׻�\����!�,|�����>��;�4P�����C ��������!��Υ���x����aՊx�����w��`J<�z8R6.(О�ϴ����)��g�2
���u֊[ۿ;��>���	K�k[f�PKlc�@c�S�B��~�YBX�S� �˨Y�.#ͥ��Eu_\��=�\]�$�a?.@�����-oq&JD�5��ϼc�O��͊�N�t�����A �li��?��s$��_Tn�T��R"��q�( ��nI��R��AM?�0����{���gh�vq��ϛ��œ�G��c��\A}�'�؜�x��TCSC���=�$�}�.}v]��5��A}�``�i�I��U�n���N��bi�s"7�&p�n�G���Aq8��hi�I���0`tPI/��׭�[�ލ�s1�P�#����������\4�.�A�Um����z�yO<,&�0��sEQ��C�h��dH$��=��P%`N/>JJ�	������t�)F���j@���4<�{mw_�0jM��r�I�W�H��!�Q�D�v����e�
�v�����{��[�Q*G.t�ƾ#x��ND㷂�U�1HȲ;�����ĀrL��a�� �w ~I�6����v�*Bn�|
��>�Ϧj�4a*�jo!��f��}Ck�oﱣ�n����*��=^t혧R�BGFZGwu���;\j6��MA�8�)�L�|�ࡓs��wx�C΄o���?��%]e�^x_T�� �$,��X�(��bs��ש���i�������So��	���.���)�H	9�2��7O~��c��U2ʤڶz:�I�ϩ���3^!:Os���q���D�s���%���A`�Į�BY&�Dޝ����
-�ͣ!=�� �A��;�f��k3@��(�N���Lv��K·}��ӴV��*��IU��Z'"��0����G �k�����4�:��E秡�N�0���F��5�_�:��{ �ܽ�k�����J������~gS�l�����
�P����*�T4F���u��H!��L"�I[ER1����3�t���[�>OB��R!ivx�4k7?���(����9���,�)X�	v���T$�#yE��G�Y��H�)��Yc�eMtFy�<���(�H��߮�~��C���8�	18�0��E��_���X�a����4j�ݡ �iM���=�:h8~���n���o���F��ܵwRx;�NJ�Zt�΢��R��Yz%3o��bI�0-����|!S�u턜�9^�sq����1ӼN���q�?[hjY�
�ęV<�9���Gn�I�V`=x#a%N?V]I��p� �9�E���@�^�P�>�!_��>�!+�����u���´��yJ#U���Capx�a�1_�D��?^} �!�5׭ (Zu����
����(��I��PS*`�;���<g�r�D�(6U��Z�Je�[	�B��c)��\7�r�砵��a{씈�R5%����M�q�&J	o^�iM���p0�5�w���fQ/C:��xpYG��gN(��5�Q�B2�"~D�}��p]�+�Ê���C��8��1�1�,�Ai�%V@��s��Hp!`G��8(�ʾ��e�W��)���sZ{�<�Z�t)=��ȉ6��j�c|���?`���)�U��3̏I}�߁`����nU�O���{��N�q� "�OHj ��g�Q�����=<!a�K ��vȉ�=����(��P�T�2���)�Z�'9�hЯ�^��sR���G�	=���h@p�m��)5�.ȯ����j9����{���A@���h��i�f��E��?媲��5�j�B��Cګ��d4\�5 ����R]����\�?�9"�H�F~m����,�e�
���v�J�!�����7.{�DU��h<����u,G5�u��R�����;J��?AIP���-�"+����O�\�Q��#!l4���)��F���j� �8��s��ݧ�s/
�"�!�|څ�PS��~�M�"�I��(��:&u���EMG>�u��RoPe�����cP��Y�����T����o���9!3�S��S_%+��0	7Hk�H(��7 H���B6dr�h�#y��_�d_KE�Aw��w��9S_�4�\+����J���Vdc8�?>��s��	:VX��'ߊ7JP]?���T�l�mmpK6���:�=��#8'-��fۧ�(�Q��>�!�[���k=K%���Q����N���bמ�$��5��u���4�9�Y��U'���^���U��傖 ��$Ә	>�V�Z޵�'�$�+�$��_�w�)}^*ҁ�1X�J't`�IY`9���d����f�X
�1�19���rP ��wdx �a�����k��­�ct�V�� 2�������!&GX�R�.��6'4ƟG⨌��3�y��ߋ��2X_��{F�#�G5��W� @�ߑ���ɎC	W�V�i��L`W�WHx���RX��@�f��[����Ჾ�m�ݙ���1�:<D�����׈#�7��9)�ێv�9'�8iН�4� ������K2q=U�<⟸��?B#�-��i����<�����8)�F�1�#눛�������1�J]�G�^0��ug�0�ɢ��,�+�<텛:���F������nXӠPZ+\���y jN�H�Zu�B19��4�y(� �C>�i���l�����Σ��	OA�du%F�>\6OtdW�/�,��˩��f�q�ݳ�5M���������m��t�jɢfc�n���|�2�%f3���;���a����AÃg��]���A �h,���.�W�ʣ�!/�U�Y�"��b#Z���^���,u@���@�NPY��zma�O����/�<O`b�sH'P#�q:E�u���U��F#��K��Dtqܰ�5�O�%
a>��p�}�s��L>d��	���{_�:V�Z��T���-\a4��}�Nz|�t�k�I>m������/��}��6��Q�B�y��5��7J��%j�(��M�Ql�U/ğ�`���gI�䴿�e;&S�����\�����^u�CN��	P6���JW�S"�o��4]�O>��A���bD(%�^�P\9?���L�+��k�����VG��tMm�8[�g�&����M&����ˀ$v�J�$����߀	H�z���._��Br�x��F��-R��%5��9�K�G�����ך���խ��w�)!�u㋟g+��hb@XfHb�w)�~<?�����^�:��3�sAxZu����]c�˵=@ ��)#��,#�%6=b��(�]�"�4-.�aPؽ��Y�;ZL����f~5��ý�a��hP3�t_�F����w�I��u����T�� �i�
���ps(�oZ)���t��q۬�A��追m�cki[�h�j�uJ��;�:�nO���
:��'pH��W;�;�M�Z0�35m�.n<0k%c�^�e�Rc�;H�=?׿��!��E� 6l�͖q�6�����M�7�f������l��Y��rS=J�@����)�-~�6���N�<��'L�&�Hͧ@�$��k�/�o��QR5e%� ]���5v�t ���'����av,�}\�Iq��D�<]��34��O-���)�ԛ�^�7��|/#��W��[��4��l"���w�AA;����+���מ־q�v��
͈v.~��Lrz�Z���g�n��ܴ��+QƂ̿<������\�9I��b.p8`�؍�s�5�
6Ƿ��XH��R�-�l<���u��j�zWW�$&.ё�"�_А×�Jߟ��.�]���"��t6)6����!��P`C)�G���$�hp���P���u�&7+��'�f�(�4��|�A�r}!��t��~��s�<�Q���פ������m���Ve�q^ ��)Ok��	��ɭ̒��̋~�*;�`��8ۓv��`W� Ō.���Gq��V'p��S����?y�V~Z[�PG<� ��æ"�?��+{�<*]���:���2�Or�H���ͨ���"����w�Fc����a��CH����缽����2R���¡��ǹEUr�&�c<��N���R��s��yIЈ��6%�l�N��ό��:Y���/R	��\���.�t�D\6���:�����S���L���f	��r=aO~x,	��W�������s/E�R��BPl%�0�)����Ԣ��I���T�/����R�8��Mx�����c"w;���;�T�Wa�+�Vd�a�^I+#1"�}NX&?D� ��E�����ϧ�F����}����׎�>֨��YX^m��8X��������a�^.�l©%l�-rͱxqE5 ֲ����}�)��/]���4ϧ�A���1w�a)��nt���-����^��
b;��dW�W3w�cʀ~��]����H�?��7ϋ�^m�j��!~��寻�&]��EI�J�}�� 4�����e|��4ɂb� X=��$Ӎ���,{пrX�,�}@N��3���<�߂�:Т�X�ʂr3{��J�CD:z����jb�1:LK6�Jk�5���W�R� �S�q�b��_کd,��a��F�H����yz��.����p���#�ͫ����ֈ��ׂ§�־Ѽzٱ�wIV�	��  Ϻ�3�����9'.��Dt�^�]夜۷����|j��b��?�X'�4;"[��܍ۈ�8t�un
�����U�VS���Nz��i�V�g��o����T��2�C���Axh6�vmt�ԗvКmL`��!";�K;�h��!��-$���l#��R�yʿ���);�3�`<'�ZH`�i�t���v%�gd��Z�ǫ-&��џq�e���x�m5JƳT�b��T����a�J�+Í�UR�	�{5��W褁LN�=�'�<FXyP��[9�7��u�.�����v*�al�S�2��"N^��wa�ӯpNcG|�_cd�3_B� �jNڋ���ҧ�	`y����K���:��2��r4'�}���gŀ��7�]�3�.q�-#	�:r���JrAݿ�I8�ˉň>Ԯ�}��/�B�q�P��ޖ�`��R;�Q��&��M�\�dg��w���;�!l��t�5w�e�zK�M��e�7��݅�4���~�3��v�m/�<�y���ㅙR��"��"(��V�ki�!�?��f]סc��m��0��*��t�T�^�/���Kf��?����:��Ft55���@h!���j1y����$��o9X]9m��k���n�5��į�+���C�Bm�n��48���:*��g��铜���������J>W�	�׎�t��-qq͗oԈ�aW�L�G&���;�r�oX�AU$.k�9�g���0N�����pTF�d%�6��M˛C+��?�d�?���j(+z���e��sE2�����?$����m�s¡&�'��WQ�.�Jq�{����mX*�/֏xY���r���M�+j,�1ض�3�`�ty^�ԯ��n2�O���?�<��<���ܧd�E1�ߨeZ)��p1���߿��ef�uSL��9:��:�T�3!&ς��al���L��m�˜m�"�T�3���H�5�u*9ؤ�m�)z�%N�ނ��N�ӏ����%+�YwaKptI��w�	���Kxjѹ�z/�;�\���M����8�]�vU`���~�B�"o4���I�fL[F~e>^�z��%����Jt���L���sZ�=`������N��N��J.��E�ޥ������?Z$5+��\�8��Ou�>� "��^ş����諈��?Һ[&7*�Ti����"0������e�f� lP[�@�j��!b����Z�	Bc8E3�7RpF���4��i 1��	ZW���A3n��Q��X]g��@�I��M���� 1$!5���*��ӣT������L�+�=2T�qY����e�h���ef闾��Dl9�"�xHŒƞ��N�����Ha�V�Ȕ0_��tv��B^�0��-�=��RG���Zb�n��X�$�<��j���Rޔ6]׸������i�b��Y�U�x�b�>v-�U君�}�\�:k˰`\�d��k�-����<~�8������"h��L_9(�-L�1�V��
A��K�V�s��e�\+�v->6�9y���H�׬�(�#0�~�G����}��`?@Q�s�B�"��Wpŧ�OΏ�g�f�<V�O���U�xYXL�2�(9�T��U�P��r�-E+f�#ȭ-(��fM�u�~8C���S��P(CZ����Vs�B�_/x����h
��:L��"k��V��s�ı)������J���MȢH\�ջ`Q�R���ք,�U���P++n�t��DU�����g��gG�[B����U��ֳXs-�,zqj?��&��Ɲ��0�3���k�튐9��D�V�q�a��YW� |��ٳH��J�"&̤����$�OE�o��z��{'kI���ː��7�C'E�m���Cǭ}y㶍��R������ጥJve�jS�Iu��%�e׀�0����L�Ӏ�@.�N���H��Sյ���aT��}��{����X���ث7��?��!��Ybg���}�����ZsҦ��rΈ=9/sj@���7���UC�M[�,��͟
�.|�E�'��j�7x�kH2����Q]�ҽd��pPd���/|����Xb�ӑK�\::"������C�/>��vk�>���;�R�-�?N\��Qm��3 Ĥ����kO|�P��.$�/Qq��2�
I�ج�?��(�.�D� 9�2FΈ�vT��̬G�2���qcb���q8������0�w%��� oY���n����m���n�.���[H@�x�<��8F�\���
M��g`W��󄧊J��RE��s�"k���w{�.�9�Hߕ隣N.8���!�}�3�
\��@�~�1!K�B�n�����[azI>� [+Nj�?Q =%֜�y����ҤIHl��R��� ��U��ƅ9�Aet&
��P�-���B1��#堦��A��ȷF�ק˵���EM��?���������l4����'�KE �s(G��Q6?B��	�^�sW��Bp{|�|v���*i&��]d�]�-�j�o�_Oq���s���sq�(��t.P%�{\u�NWE�|=ꖦ;S󖁻ˆL�d��-nX�g�O뺩�-~9��J�bp,� ǜ�h���n�/�05ȸԘF�X#M�����g?!��;��f�'_{��N�sCi��q�����|�g;+~�匍�:��_|�[l���l���b�V#��(bD�~�Y�^yC��m����IM���Y�ƙl�`�l��l������6o��KD �|�0OWR���
�A���H/�e�p�4.RYU�gW���q;���Y���� G$�&���J�dE�Q���\���@R{z��K_pVUh�8�?��[oq�gl�h)�N�^-�yI�5	tUo8X>��i^qʬ������{�4`ө��˶��ۑ�])�^D��~E6�iT�jBj�x?4�ѩT��D�<��&^���vzD�4�~�5�JI}��#M�f�N�~ĉ�;&[�tw�����,	��䲛���(���X@��N0c-4:�S=&W]�6�`�b�K�!*M߲1,d��n\����M�(pRR_<�C H�Iw�b1�T�c^2,�c�����MxP0'�)�(ըM�Q��[̍�U-�>=�x��� ٵ#@�U5ԴF�4��au(�݇�5M}j3���e�Bil6p���Px�l�j������I0c9G�V��l"��&�+�c�V�*{�?ZǸ���@�b��)��k;��NѮs�����A1W��=8t�
�q���}��
�<��^P$@�#Ҕ��N�؊��0S��(+�H�oC]��"�_�e.�t`v&c�M�=e@`�ch9ܷe_�\V��uqvX�vE@k0��]�Lq���^���#�i��PH�2%��n��*C�(��\92c�F��ҝuI��vA/�a�%i?TZ�6 <y��8~xzDz��X�IC�t� ��1�r
]��P���M]�r02��g{�ʱ�-Gix`����i�v�6�E�?��L[������R�arZ9����xM��?��]W�3W��j,R�4C�gq�}�ןAR��me8�V�>�Z�d��]kGp��=���2�!�8Z0�*�����Y�Ӆ��2��X4��z���S���4�g~
sR@㐓2_-o��kg��`���o4�	��Q�$	��8��O/��R	�x)f��.��ܓ��^����-O��@+5������Y'�+��T����#�X�gE��ui����Okq-��!hth��}���n��Rl>$=-g�궘ԃ�	L��6�_$Kɧ�.~V!F.-�O��
^�+��Aq���P�:����:xc������/J�����!�T_G����U�j�'դq�\�uJ��u\�,]�1�[ñ;+c����A�В�7|�
�{٨ˈ�-U�YT��Y#�-$�K������5�qe�?�G|���n],�u�I�NN�jY}��<1�w �����!��m�3Õ�W�Q� �,�� Z��� ���k��"�$�+�5���5i�K!a�*Ԣ@��Y�|ZKJ�&+����x�4}냰_�����g�^����n5����ҳ��!�*8�Y��*�jݛDS�I��22[�����PNlLn�ʠ��var�r�ws����D�G�=h���![�7�Sn�'�%A�CR�ɩ�k&[5�y�����
�
�$�
1?m��(Ӡ_}R��bz�-5Q�C�i����J
t^<az�xw�f*�?���k����<�m�a�,(���1q[QfH��Ț��y'�@�U�o
L6f�Dpv7�mZ0ł�/³�s�M@M�Qҳ�{,�5񲯮����Yv�`���@�`��/<#�4��Sަ�f�n��i�Ϣ���o���.({~-aG�<O���`ŧ�,�DC5�T-%/��c��#��ܼ�΂�9��%?�e3�HB�t��K~�z&�H'NN.J\��;�1�dD+�	�q�=�	N�Q�%
��b����tp�@yic�O�Zr���T�J>���/gz�*�d>��ۭ�]��-�&0N�0�
HS4�r�		E��]���ψR�$^s^Y�]_���ڕ"��|��y��X�YI��t2E�gi�����a��7 �%wg�% zY�����℧�z΄�P?�ӹ��z�6�xl����T�~��J��x����Q�	�.>H�!�X�>^.oa���P��	�j/�tV�2E>��1��r��w/���<�>� \���I����@ǋ���P��)2�[�ki��MH���u�Ż�����el��6�(O�� [@����ّq/��&`I�¼�s��鏒{C�&���HU�Z�K%��m�5͎!�v�¼��yfX�Vi����J�[+xo�z��X�"dn����}�ڟ�i���ā:ܓ�ғ8R�q�j��1�l凩����ԑa��Gg�B��&�x�)(%ӯ���>��'�ю��5ҒX|��|�N^̱�f��D#p�޹����*��ɲ'm���=7q]��.p1Ӓ�Z��q�&G��
H���٪���΁x�Ĥ����Ǐ���Y8��up��g5q��[iN�K��T������4T%�y����\��.��SD�7��;R�����vu��O� ACh��zA��Ugu
5w҇��a������#����_�>��o�9_�ɫ�&��};b�A�E�d�C�1�@Rf>�1�p���u��}qNZ���Yx V!��v��A� �nd�Ĩ��&h*����ؐ�����<EŮ��m:$�oG����<�sND]����Cf/Ņ�4�!�Ogn���!��� ���<^���q��G-�F"��1��|���LL�O6AFnH�I�� ^�m�y���v���v�Ĉ�Ҍy��fq��u����.��S�_�i6���i�}t%��p��9�*����x���Vh�r��1����	IP ���^�uA�-w2TY
4��cyM��4�Yd�"�s��u�b���v�T��ά�3U	�U�w�R����ѩ�/�J	�J.��@H�d|��SC�54�(�%�s�ȍ��o�+z��H���21����?1SCI>Al��1)W���Hì�*i-�VZ��甜M���a��	�M��VS����]�X��u	3���f��:c�#�E����پ���q�Щ'NӺ�_��nr�)��\���O�}R���x8�A��ݨ�4�滰���E4>��8�`K�! 9����g�z���홂 y_Qp~���_w���t�b`Et�u'Jw�E7��LB�-r~[c�{�Wf/�Z.T~�M9�_�����Ctו�N��$̜�����蓬:�s��Q���?Q�?(�ך&�h�*�e���A?d��Ps����5��U����Ӹ��������7
�����R��)���@I n[��Qw�J]+��7��h�C0�k�&�;~��:�Ui����-��r�$m�qη
�,�Я�~��	c˙�CY�?��B* Ũ�9<�	�"��s8�Uwb'�8�.�����%*4K���c(@����U�F��*@I`(p����;�� ���B�>D0�;wK�UJ��jp^�K�0�D�˄�m!xU��}JKā2>V������ev唪ٵ:���zk��5~$i�v�/�T�Fƛ�h4���p�#��c�~.���E�"c��%vt�-_�F�Z�I�t&����C�x1�g�͠�m�B�Hj��f�)r�螃�s d�b)oy�WG$�B�;Z�?���:)� �Uo�o��E��)� �z�UZ�<ż��f�	�d��N6 uK�.M�D۶�,w��n�P3%8�(}����]�X�]B8J|&�x����|3�vGc#�U� hsG��:`�
���b1�?9�=2��$i��b���ypwoC���{��>�T؎�!�:C�smB��[��+���7�@�ѱs��'�ң;�����^$��/���^;���=�SZ�D�Ƭ`�z\��U݆YG�-H��;�B+�����$����8�h���on��OlJ#J�&dq1�3j^<���v��ٗ� �G��!eM�
�_| @��������v��=���tؼ�Q������=y��3��t
)$�V����9�3����(fz�I�� �V�1z^N�bK�<$/���1�Ϲ��v�� ������F���n9��>p��J�#E��\�x��ؼ�0�#����E{DFt��ݸ"�K�̱~7�F��*/��:<_�of��(�FB¨{�)�����Y�Uqm.�Ի�G��dW�ٸ�N-��־lh'in���F��iBpЇ��ZT���h�G�	2u���G(.a���?�5j�v�s������H�3#!�~aQ��q)^��W5Ɵ�*dY�ؽ����W5�ص�d�.p�'�q}��<���ZC����ha}�� |c}��C��O	���m3˛,�����
�Żt^AHI<ڝ��E�n��.:�~T�����(�M�"�7)�(A�>�jfs���7M���$Q�~k��NkGxn�K<F{���j��M���|�m���ƛ�[[֍�N�uP)��2R%@X�!g������g���*�u|�y���$�i��"�"�BΌ���[�
4H�f��f�R��4�`�v/��rm�C~���=�-�>��~7����Yl�<hD�c�����_9ޟ�c��5�D�kk�)���x�{�Hn�vl��#h7�G�'&�.5#�Y�=d���F��	+��iJ����d�a��Y���#.���8w13�EA������Eu��z�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               conectix             1�qemu  Wi2k     `      `     ����u�M���<���                                                                                                                                                                                                                                                                                                                                                                                                                                            